// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UtwDRyONbmIhqB/dD/JXWx4aD8DgzExkMdReXWCQv6C860hLr+FWvaRM8NW8
RawEqjK6BqaLlXoMksOwYuAMYfN2qXO4cZEHzV5i6lWlwIbC3iIBUyRHv1wc
Xs/bI9aG2wad5g8kYteNFICbD4BaQ14Szvvipk5FSNui9R514EDA6UnfJjrN
sVJKDFR0ADawqr+iHgkfO5OYBXvPdOuQLhQMobACntwv+7ao3Vw/PUzqGbaM
NRWRSlLz7ujyvBJVLO+atXR1ojw1UZkSiZb3HDt6zK57CcqMNeEsvtFcY1pa
gg4QrSyoaL2rd/s1sZsaXvwLay3KGlKgzhMcUCNKaQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LHMCXeejoan/dzHSnvssRLd2S2FxYwqnU6Njxps+0F9XXTN6ZFhk4j8xAsoG
UpOZGW+yXWTbuXlj1eE8ubpO6jS/qBeSusiueQGHJhR9kHGqrAHEAnRo2AwD
s+0f0yR+pjfw0ebd/l0cVPJPxNlMob5qCxQ9nPVNCAvF3MqEM1r6UVCTTYfD
sF7pbhCZ1WSEMxN9Opag6vDMpZ/RgpbdRJCDnSiNdVDbraLS1WtbLpBkSZj7
nhtiTkjKwZJNSoAKZO5A6c0hdpN9fUoT3A+JAsSdEuWuraHtHBqIWwaQ6L6g
FDxtXvz39hc8Jv8MTXHXwOPh7KhqUIwj2bEhq4aVIQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QgO477kZwHSlMqzbMVxUc3P7zJ4Uy9NSD6HrM22SOlu35427JnIGPji3gAlK
4UKPvP9VEGgd3GN2lDhZCx+K0cqNJQDI8e9WSkFbcGuQbGOmepDkm4oPZawY
0mNIVWflyKhrsKrZq/wqirya3sFvqtAf0b8p9fYfGIeITYZzeVT8P5dMRjnB
inXPmsRGqadkT+M/5WkuXYhr0JLrFiqVZSFGu3FsPnsdhw3318Ixhsd0SBHS
+t2fJvfMoOZ45VS6htFfBa+z2H+z19/QCruao0U9vZWyDMMzq/Fx5t7tyQBR
rHlGx79DEijfDrG9kBaEQpjUExxuZ05MC1g7oCFfnw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rd+mJpt2n62jTEq9SPYuP0C0x1HxYQOV0VqoLY9krZuX/3epsjt0nJCk/axX
akLiBtJVQM/wPcUKftV0sQPD3eGjQxFrGsxuYE7OIwIy6Oiq29WVd76b5aUk
VJdfqvSBqVevKv+pnSEZTD96zP/AOSHSe0iRxgNZQLp9mIhXCvk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
prOf/9KTCZfMYz3yJ0U5xl/VYpBjmkRLTLaszYT3ND42Fgl5XbTor+NiTG+n
CXb0cDQyr+CPbpDz9lNHR2H7+3ME4zxh6DGk9n0P6Y+ntjJEj/bNnOZmYeb+
3PiAztTwQpaNGbkq4mNRxxIk3I/6Gy7LwWthOak4SmueLbct3CNsBSgkqQvM
iddyfgPB63oeR8s/2vjWpwzCRwM+CXMgv4nSu79aUsunbPEET7jMiKDvomhK
W3pRfEIcpMxJ+260y7clNRbygYa9fECgNbri5LRLCcxB033kiHuuY+eF0pJa
OOQY0BN22SO4Dyxg0vdt0vAnaFqRlbth3hcGRRJNe9JSZ3gaKF/7ifkn3Ni8
A2yy65mowyox6sCf0EUbfjCEkKs+SeLLJ72LUpz5CQuOGuFg3Q5jTMLSc8kP
rMndr+IJylNBOmsvVvewVh/DLu2HCS0sSNeT//5S3kE0c6Fux2uPWsYYsIMd
asP4ezE4vbedGtVH5QODCK97Nv3+eSYt


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
F3kQQfVS1ng4grkdaeCwM3nqM+CQ5R+ySR0w3QpfwUkMUGL9iXOO0zRi/u/z
NGH4usj5L7nhcchK4fnoLrogPwz9QQ12zgOrmdlr/ewobjRH7apgPrfhySlg
y5nMMiW59r52wnuUKtq4QtJsdU2Qewtp36V1/4GLrY3QIDAQbOk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GE4jWCeuHBG6SC5zWaMx0zmkXBAAQJKVwa/Y/H5ck20S+kWYUc0C3dUbWZfa
KkY2rQITqhe7ZhBQG1IAIUcQQUKvoqvMZ5sYWb7iN082W3Dz7JruwP1mqF6K
mVDVZcK/mABJmg24We8Dkp506SLcW+thOjp9/GxLYkpF3qkhqiM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 18912)
`pragma protect data_block
ASiv617W59WS6a2uuZD+Q3ujSrCgTxbO3/oiOAQl44UuzJ1YwtaZ6IBlXBST
3Rs4uk/nj3rXNSNUSXZj450z6g4e8sG98YDIBOLxnzVATQYjIjacKOdj4SZN
o69q3JFnDRqGpT2UQaFMGKmebRjfGyZ81Dq3R0dnZhVs9zWyr3xvF5XZturb
+mb+VVgE+5ZlZMCq5bm2drxVTBuQPMI1UvAGmO39YV3S5H7kNAxzfp8/tGaJ
YBu+UDLxHvxZMDUc0ovBJLMkfSP4peXFPCVUR7nVEeHR0XtkblP4XSWAL7Qa
hw8FJ97Z0sKl3ixrbiGJD3Oub1hrEzRwCgAP74phTEvriX/n1UK9WoqfbV03
JoO8fTr3ro+pv2D0ji3ex4bLDumpHxwginUSTRTw8QqwAoisFmGjc16dDD6h
UbDX8PPDg0J/QfcZtaRUXsB1U/I/cAlhpn6VaiiS/AZ66MvgD7xc7GWhwaC7
hrPvkfCALogrmgFVfa3CaThVPQxXNYhGzbWuhvGbKFJCD2Uc/6nL4F86voWe
Q8R16EcCpsgh/YgpEKAJsSwQEEIanzXDAdkBy0Ztq4rVInXMkLwBluKGkbz8
Uor/ealQMG90olTuQU8tXKP0gR+FiALnwDb4xohu0gCuf9ZutTMy2NMnUUwX
2wNBflSc6nvmCd/FAJSXtuxL2Nca12hqn4dgeNi2uf3KrIaLREuCGD2iKaWU
DY8PYKx4XUzdfpq1iYVVcDnj1dZ+bnjfmdb5Z1W1r2c5uUl4ixIMTL5qGaIW
OHhYGOxHjYvnVV0pIDqonQXOUptxDdGPcl4K4PADE625W1aujJD8kwvg4org
Mq+9E9DuddPrQx9mUX4iNW1qN7SJjH6etDo/LLKalq1VZ4SDxoP5AfzKEGPt
8woxvx4L10jGZDE2NGQqsEEToQs51aZvErvLFgssVMCT9zU5fPYlzZcT+ZH7
XXrUBqoLZCrwCCNBhEK7ru/DVr92XkZSaRyXq8a0ohs+ZSTecfiP1mfjAzig
0SGANpWXrJxsgHPWsv064Rw67GB05l/NJmWjqGK3xszd68dpgPoVRD8yDDmC
nH7tGaJ9ciNjJ5bRwV1/scAATF/tB8sLxMHIunSSDwL21TDGMDjnKwecRkg7
IVJMsOVvujRzwga4dmEeaDrj0eVKR246ZvsVlIffQjsiotMk/KfCBXaUSF17
yY8dvv9ul6oy5ESBxuFD7PnfVL9t72se7ZxMVUHGmbBdP90Sigx2I7LpxYdH
+/yeNLy4ic6IUYrTiI3qgssa1CEr/XDJq4l2Bdu/45iQT5heQi0LMhbvVBaG
9rJtAW1LkTec7UVIZTiFaBXp+qIAqH131h5qjZQsy9iOBYNC2My8R2CBQnn5
uMcI9h12258id+06+Vtb0OVYD7wsSk22UqXtcbpSP6rb6uTHQPR+8w1vH12s
pXvLMt8t1wfnFp+Syk2ckMMeyxb/Y9/dEzhnzqB1VLwETAF5qwdr4PShtPXz
cZNUbwedGia0qxp5ii/XkNyTqwEBd5B/ZBJ8q2iEwO104Woo462QY2geiM5u
wE4NJCOBIpG/J3OXV6ghjcTA9VTz7x04zpZsLO26EWZKbfXVABd8H3MqqNoj
/zy0eFvzqUsMYkIjdw6f1acB1lOxvhUVP/XjN56Q+nRBeOkmbCstQHClm6x/
rnK5vGftg4IOxZvLW9wxchiqWx0DcEGVLzJXAmBVRWfVURBQkM6WMHvupagh
QagQNlgH0w6LbjEI1egFsD/XygSk341I2lgQGrO1wH3L6DirzE0BquVYZmZ0
rFVxr05LRCBq7NG7XyDRoPQqM+XUFBEp0cKLgkXQR/JVAWpimF0pjld4dh73
C7tEd60Lj54vvI6X9EGct6kKb6gbDiJYiJXVUdazVAR7ys0G4zY032FdpuNm
PYqCEKTlP3pKyp7ktaLCYoEf01DVxFdZD42iE/gDdouewEXfXatEpZAu5sJX
2CNs9g79q8MW+N8FDy5UtPpINkav/RTaR9f5eZbv+B1ymvNsuiDERFKqv5VX
DVg7UZfs0l5yjPt3H4htIvFBk3+cMb4e3GWANIkt2Yfi2UcO0QthFwBWrb5q
XZe1fC6krEt5y21wbYpvuDr1/sFJ+8rjX3HNtW1HbCvbZMgVeuZGs+1oEq6D
3GmNfjeWDkD9LQE5xnXfnb5OmQPNVmAjQ6gUKA3MUzGnEhhZ1UvTOCglU9+h
3Y+Fv2GKTmFdvIhYeYX0jUKJ2cRah3dUYNViH/YHSCjv6tiUCMQUE/UM/7JX
L7iS2NnkBRm2vmbhMFActu6JjDS4gBhIozQL/q8KI3mK37x8Ct1hCeqzMEsx
0kKf3m3jTnypLIfuoE13E4JTvZRNyo8Zd1BM7gaB4DM3J7IbaPPqnXkxLFT3
Eg3+HWhov6ppGrSGWaZNBqDf/qcqkl2GlCFt0TGRpaqSBHWV5F5co3ULROiA
NU+1H+JN1NC++RzQf5xJM65gVrUwGnL9cLdTk8gRANNyo0I2Kzd4TvvoCaj/
KPeJI/JNDa7NufYmE0x5FHdBcPfC74kI+1y0cMPvUXP5X/8GPdOyHR0+/clU
V2GQQ6otXQWRkCfP9kjhfTubbqeEZMD+/njJfGXd6CzH9GCQTGDrgmATHA5h
sWk0Flm0aYQQ1U3hXsdivEg1LSWca41CdiCJGXU3MotaQtwX3m3gyVs26wn/
B+IUDhxwA1HnhejOLA81jymKfClz9HgPcU4CQNdbc7KulMYReNIbYbAPfpYG
zOReFAsWgchZI2qEzuJ2jgYsS0aMuj/rJkuQDOzSDpn5JQam7rwepNHIJU4Y
jwfAaj8Bd+2Jn/Ohpzs46mrqkiWBMx9b9hp+APOYmQR0EK+i53Kptl7QztAc
nKppBmHIFrJjriKfiEkCnmhhWm+L4kG2++EMUPXX2wZQjF94Fg35j8MR3/kW
tXL+VyzGXoGtdaMtUyllSDXmUcQkqlhzE9rhaZrejhNNQSrP8iLFuauUrbLk
OAChrfMyfK6cWNcfJM9VAxRYA4S9QfPMosZAKx5IrZ5Rd77CWRKviOEPrwF9
dY3FzUyzzeGaMwjUL6+FEOuaLicLQ0FMC4SpQo9KQyu9BpGnPI1dFU2ZOQVF
LkoIN9mMSv5qqosSasFTDAl3anTw3sqih0S9jSdj2e+LYFzJhLi25McD6rdF
nEklL/IjZXX6IpBk8VNbN8sHLlEapEkb4m8jDvcZqqTLFM6PSdiZjEgWdW4p
lcDiXQhZIhe0rNv4q/OwMInbyjScv/xnXEw0+TfDBXcswXXN94rc1Tn1m19Q
ujKe8MxHUWSoRLj/9j+CPvTVvCWi7J1s7HQ6Y9Sc+aatsDTdNjJyTXbBVzr+
ae2/xNQ5ixyuQnLn0ofYOjS2KGjvExJUh3a5xum+f/WNICSeBk2VhnUGFN1v
w5PfULbiEpFV64BKu3z+BLFwF04hPcyI+uj34fLJBYF/11DFHbLfqXallhTE
QNS4sX2AOLKaRmqVdS1RCdMb+Z0IXU/NWk2W96YRTDIyLsUR4YO4dbBde3lb
Yvr5eEO7ET1voEm5RVbzkg3CwzQk023VU8WBBouZ1hch6LnRzQuJwVRsHz04
E3y41t1meHUZWqJsMJ7AFQ9TEiKwSMaesZ+dzfwr8UW9ir6qC+51JgyvQmtj
2xh/CQI7hEilQiKKzxEaVQa6Ptc5XEd5jiNN9UuXb//ijAXLWo94MFPbFCVW
KczLX9Pd0n+jNxlsRVZeoigHQGEAfRYDZQ6tkiJ+3BJ4Ly/Btun1S2FXdC79
9itWR9VCokFae/3JTsg0rKukpS+Q4A9FCjbCBB8I+6YGHVazZv+pOU6plN+n
lgmkVSa3QwyZGlN6Cu9ZpUVqhT7vuecvN4S0jrcgIpmSxkkM/eBB8Lav46MJ
EuLtuzSGpc7O5WWuFrMRrVRGXBh21IcYJfabNhLFISfAr7nGpeYSXOVQtQfi
FgxY+c2qWSeTZYouBrxumNtuVtcxTXCxDmvTedwbqSblVOO8rPnhngPlsSvz
zXRU1SEz4xzRa+oL5AwG89J1J1G8uzs6+SW21VdMUKkPeOZcXj/tEDwg/y3j
K/c9hVaBOCXuvpZc7IJg9t6sh8UIj8DferouxvHomTPY0tuCm5mErmhKyMW8
Zs+MiMKdRp+I04Yr2Y7kkbjkqI/n28ag4IaIWCp/pM8R8rjIFS+e0LvogCYe
1HQu+wgv0no9qwsOdbKKCOVgMB7wP7Bpb5BZeFw2wRaa3/5DPvXalMvjeldd
0KngIQYAGqdPfZl3bOOFWfrbU4OhF6Dr84QmOYjlLhQMh16h/hMawpbpKSq9
aapCaz4hq847y9wDypIaAOjKNX9J7tVsmQzP8EMsJujd1Saew3JyjifC2XD2
En47v+pkYSPww/gRFEGe5UAg98PBgALhGUKkIXLsNlpgbfcf7B8dz0J8PjVV
pNEwwzFgIctUHBLHCD8GlRiapZLjn6Ct17wFyZ0uZOrH66fhFpX9q7K+mx3x
XEKFoj6gzbahqcsuta/x3y0wAxTzDedoJiMlCb70Koae/FbmGMwA+6UsbJHO
+A6QJ/eW9KlctbsDk9hopa98/5H+Mx4WCKBzH7uJkiP1tFVCCfr4Fdezk6ON
qmlDBvb8PK5BzZyH6GaoZ8wk4UeCJcsylqDXoyVPEekHLzcO96CGJcRDzT/O
m/LpuqDmKw4qTzwWBu/yftbffFNIu8hufNjmu+hsfHSERclfCI75uSsos8Dl
wbqLNEBO+aGVv6tODZDbb8jnAvQCWHHyRw3V2YTLKdLs06tkdNkVmqelA57v
7HfcdLByAFzozA5hvRdjpBJb0Ug+gN+PO86MB7nZC3HAb0jXFhrSOkiNKYwS
PNogMv7CHr5nUTgJN/WHO/ZUM2KgbDTcNAt9VGilmOV9QnC1gDS3zj4OADv4
yMyRcXclOTOgdgbDXgKzW69XoUy4pkYAPNZhRw8t9sJ3WW+ptITtjBbq2Zxy
IQiLMEUD1ttNixlSUtKCH86CHtWAMyTN1aYmYqCzSIR6vljFALIU/uuTaiOj
sWzznYe6N1N40t43DI/F2D76ZdhYp9lMSyb3+mN0mJPn9LG5Pai4Torp3yPa
tFRd0nSl80QuE8T/tf1Td84siA5wmwDWTwkEy2il4+z1iX9UCLq8KR4paiyn
md0PP8f5snzyhz9Vu1alsYv+Ch8c91uR1E0RyBH8zo4uXfcMCdvitywA18lJ
m4Uw2yDUc4iXRX1TS3I/QRJ0LSz4aaHvhLZ6rvKLjzZiv9XAFT3jl30PEZos
mx76a6P7dMkn7QtuIuAWftAdasEUntYOVmNCh96FHLvJ9VHrbOfQhP3oqi2E
pvJVB1FX/EIi++RqxP2fco8ABsBaVp3ttYH4Y25NX10SFElYPX5jMpHx6wRI
GUpbo2LWSpmSmDuggDf6jd6Tohp/ZRrvZuP4DUwNZ8CIpv8GZaslXgrjQuvs
CFHen80HhWS5tMMRMU31y2S098QuvGo+iBz31uzChV60gCYeXKq8Yd84KaO8
YkcB5W8za8WSUQlhBAQSgvtCSDX4huiyqWVch5BoqTRRdtHoFBAIuxPrC2lF
uf2m6v2sCyFoI0fQJJ+4Dpz4wky6dklpSjY/Wlsru03zsavidn+iMNuYOIXO
y3P9/lHZqWC64goR+89bX5o93CMHvtqsrff1umGi3zyuxV+4B9NTyY8TPkEv
QltPHrGenOgHwm3uTxFw6qrV0dGMq8fVD2czoUIT2MVq/blcApyQeD8x+dCK
b+QwFV7BLu+aDNJ3kQC3SzD0yKG+S6eQGYkrBQoedg+B9O9Jn0OvdWxYzxll
w/Ka6FrH8pvzr/ZtIO3DgW9VQ05w0J9f1BIbOKyyvTeiRUWvopz+L+BEJv2n
VHXdtcw/UQVpxXB7zUIXzZ/7ljUynL7PnTwsX+mN5uzH0Qd2CldGCvJIxwRp
ZBAONKbrgA9oWhXZ6xu1doAND0753Tl2goJuUE4A2AYBnfj6xn2Tf/v7KQ4i
BQXtob1Q94XjCeHiCBk27prpjJ8WsG5u0cswgO2Li/SbMTtyTBOLqto0rK6f
y+aT2BM0BtD1TIzfoSLt4mOh2/YxoSL8Mf6dS9TuC41pVeaaTw60RnDqiJ3+
IypxK4cQ8ZAQ0QZqXYxBDCzIT6ZFIxnt5HFc1OGxQWg8TJ4rLgDcAVJ09B42
c5dh/yt2VAq9P3LJOyF8ZXJ9d3OtnLMe5ZiCpx8d4sQBcqdgoOksIUjNFohP
+fp57dUHfh0+Qfpy5YHrmAFLNiPxT0I2qpf/GxoDeZbcJNkaYtXSPhuzr6Kw
yxK/n20WU2P0ruOpqCPzljpvQG1kh0fs3XUgRjIlaswIIg/9lgyx5ZalERo3
RRWqHZ374qODzhHoTQ9vTaCF6P86VAbmGxOwRjLqBRM2GAKYs9Sc80b94tHb
ifpjJJ8sei4bNmw/g/pADnlQhIlcMz4A/hlAvMpTmGip/h7ToCTH0pbt2s1c
s9n7XDdD/7nZgM3z95kFZluED5uru1+2W+ORh2dW+cmk4vnJQXSzfp2xg4cz
hXO4L6n2dwVucAeconZmbV63GXDxPpRf69BVU9qSoXxdiV9sMmnmWLLvKI2d
CcXo3wgsaYiNk9OAXi5FjhflDtGQZqRhXaN7wGO3dPTQSDauqJI1ea/9RrAA
RtBtSvmE4/xoE0scy5TwnFLJal12WT6fNDTfawpQ5z0gVqTPw6CoyZ0klesC
xjW0rbbYYjrNN/G0/+o/XaU88pBedV2YunjgyWMsYpOibnftt5XdkVT3hZEs
+mRIgLd97dj1NHQauno3BU10+zEa9XeRSVMMNQnH1WD+Wfxi+asLQCmNJIwN
eeKsFOh4nk2CN3/+K1DUWifDhN354pUuMz3SdYDmRhx2nKCI5kjFikY5dBQV
1jzii+tUYmjE+/8f172c89GGTnYqAjMH1g6DAbpld8STXaYmyDtTert3kVXf
XXuUJQeEnccHPL2htpE85han9TRRz1/vfql0+8Pm0VHtl8YYLKgtFFVbvAMP
I0Ot/sK4J6ljriNATvLM3O4dFYHa+UUadfwJO52mv2ddDwDPUAN4GpPzFWXK
+5v12Yv9doyeChI2mrnfI5Utw6gvKl1VvaUSUw0LFytYjvNPn0ujN0ogJWQ8
ur4NrRdwxX6eON6nmchdh6fmpbva07q5XvFjPR8aIk23QP8A+ldkblnALE0X
nGEUpwFz79yZ5H9oxWAro97MWq0xI2xs3F7HV/jTg5hoDmKrWq2iJqoa1ZyV
zjjxa35T7aovzjKhTkpM+8FYGT41lN8n7vvTuJtK3kdGeegoxaK/AsrF0YF6
PkZ/MudMEChXxIMmgj/TjiXWU7DgsBXQbDuCtYF5R3BlgKFLje0dEDZbYnBl
JJbI9dbd0IdAZM22tW2q4l1lve9OpuE2kQnjeLSkG2ASC3D6GCi2gTqUHBHM
Rwexk79v4lKTUrWKBWoQ8wnTN7nzDxHkcF6UR9aVYjlv+A/qnk8SoY38zk4K
KrNZl9SWqOx7jJ0JErv6WZN81IEnVsCG8h4N9bxXPtl5iNsAt0eaiPTu9e1Z
HitwfK+Hu7oDdYb2m5nGxUt4mXHj9qjAYWoGrzOzwRZy1Epf8EnCejn1Mwb+
MwKpB0Asa26qber7aG+HlkcXa3SJ6lK1N3XG4ozvGVeY9t4+cPr+54QJHq34
QCos5n266JKbxLWi0BQT8PrzVQB53iFUbENukKgo7ya02TJZL5VDI8cJDKbG
s5vDGDhszfE6vRCS0QQ0LAUzGVt2NPZULVEkMNIBHTt2Tj0RVACbLMk/MBka
xq1wjruCtKKKmqiGOe4dJp7E4S/5f+42AsxfePqAttJwArzQ1Y3PGPkYGgqA
Qv3PEhH2fPIS7iT0NzW48+HkstfiROKTy3tn6OiDG0qNuTwIb75UIMcy3ABA
eezWfzqA41ux56smzhZw/9OLUFYwj3PCjiHXMzCcWhyAJggWNyh3P1ZIqcd6
dXJcRVvD+Tuw9ILZ+/yz+h8YbiPb0oBnVgQPGeOMQX3FtIX0Q8IrM7n/EEId
nnEzevXCmaC+fR4ykuobfSDQNsO7FcKsBkRh2UkLjqpRHuOeBG1Z+Fv8ZLyq
Zq1Cg8B1ph9G65wXy0f4aSUxcVtYEUYmaorULtAKhwjczS5MZfTP3VLtzEnO
BmwzYQl2wY+33AbxYXR2K73yoFOtMhHLu8yMZm1BPH2DBJCF4iiJqTEIvcmn
Aldq/VAQ4u7qn2g8nMTdIsgdTsfRzwmXkBt/oZCPjcR/lgc+6RalCq8KQzul
oO3Xd9edv/ofG4dtsxzImWjiiYRWpZrZ++nEGmb3ymAAaINgMQ5smcvK0K1o
lRNkO0kcc+2QmmtN3p5z1lcVA57BNnlg/ZpjaKDS92EVxGsGSOcEmr2+L7Kz
WoGm4NXUodjNxLjp4JopousqKwmtJU770eeLLbogNDCQCTQo1qtHm7SmCLxE
KrYjBuD1GrIY3TPpzH/8jfOloM5j+iujFSnITivGYAJWv2BJuaZPg3OmkpaM
FpSn8IcxkH16YWfywRFHOJ8oFpkBahi8+PBHXQDRZ34B6UmZO/FBnSgQ/g7a
l/Bu33UVqbTtI2oUFdZO8vPzgeanghsipX1ihV/JWIUyP7W/R2gpC5fLGQ7e
ObiwcfjiXq5oDCbXHxBP6sRQM8bBpPDsLhAiyNFGui+wv4BNMxPAxJKE3LTH
1WG/GAdCWO4QciiQxUWGpArxxIcEEDuSQo8sYpXDyxS82gLnXNkhHNWA9iVe
88Hc/XzJi1qlnlkcXKj3w6bP0Q9q7l/+UvEuyAnywlJXgO5rkrKO+nRwjs/r
8FCktdNootsjRQGJ004RalrMR9O4/awLFJtGWs2gBfgUA04UyGn5wj2B3gTD
uDuYgf6NsFmfyMCdaMpLTNsZhw6vptnC2XYAAGfEQvaZoP9VcI0OUllwaWc/
FL1RGWOb+UyAGAobpp0UHup4T/licxhaAeN82p9cw168dRPWHkguHDjearj0
8GzBBZWklRZ+VJiQTTX8dI0/dnhzy2Peyg+H+emNbNRk0wmyuB29t8qrkphE
J7hY6VZ+JWCvl0NOTS1caYVa1gh4dO1Wvaap/7kUfkk+CPqjfxJwG6eJ8lRl
wp1BZuQTxmB+xo3JguRGQxSoBGNpRGreLFDIiMPhNMVDeWlIgufwbIN+CLGq
tIW1cyvq4FvldDXZlPcuhikEQZSugrtsbK0+jjwmv4hUOXSfvh/KHjQBxfzN
//KxPA6PXmQ0Wy542VxuxMk3rNOQktLueMs/z0Z+JgsGmXkGg71Y4Oo7RhIn
/TQ5x7gYaI9di9E9/j9zT7FL87/rRqm8u4oxGgIjwMLOMa75afvrxDj7fD7K
JkV56nAdqnxugs0OkQi2N1Yda+PXdQNqju5oEMq63uwaJf47W20Z4yO2dl+R
+gog/5mNQy3L19+bfNsLhoPPsRAkf0ngwyoGVYl31EAD6rT6PAJLvuYTjj84
nKJSkfta1quRa+Nmr7pZM0Ygx0tm+6YoGnp9bpw2BtTM9jmGq4ft9vzjimJL
yGdasWt3RfbGhjG+Lxo1uDLfjy2rkX8gYfhoXENEEWcx8QH9XgM+Olmc6RhJ
oJi7NJwl4oxF2S920h0LiW0Wro5/2rpnjkLpEVjBuSHHyx0mkUgRER8bfekU
shFiyQwxPrNTzEXfZB3gi2bzvgvmx+WCTzAftUfiTOn3nctJs/V/wv0xzJpq
clPzCqEENYdhwVH8f8Mt1SHtsjU381HNuNDzdJXl9DbsOH1VQ7Gvmav4RTlE
nMu5A+ydPjAyS+DjYIYgjSaS4eLd48GTWlIYsH3b6NqyD898IcTL2A53d5i4
nRjLNnpMITAVOb7x1TPrjAYrQaqVEF4X8qv/eJgVFYKYbLJVyEZ/TiHYmbqY
+D0oWyq8VzvAF9vYEyHIKabPS26iibTPEZ3PHpqw1dIISQ3qMDkpacLafcof
Y2pH/5K9Y7I8FFQb822rHiCHGZ2HwZ8yhUT5JGwXn5ZGpnO2T/3xn2Y2m2Yf
Ob8b9dUCwEZ/UNwhIxh/Ne2S4AVu2YlV1g10zMtSRy6H1C0Ga7mSyuOrVJhn
+67tcxuoM6Jos6xoVpONB45RhBL+0bMjQv9B8fmmJox0ArROj2VbR0HgzkzR
mRBrvq3XUWzCEgV3RK8iGTT1gTzQ3TzzkRl+cYdiDmVMVUPqqdcj12ghvqnh
lfg8K+jVWtgF7u577aWtxWjINjb24CpLrxKeJOPTPh+GnXcZy02+flzG+jdH
byKugtBLyo6GgvEp2wrf7bK7z/ha7OzCAdd7hiRI5w/aSg5dKGcmi9SQ/Jnr
QzcQ1zqF3X9/qqlGUz1rKGTIfbTHmdOQv7mp2UEm7RNGL0wVStbqfoKQnUWu
khDx8ZnZEMo+fL48NQxJGAloIeGPHLonFGUtOnmL5aCBrUp+ccTd3nFMI8U8
9RUfSjDT4VObMAR4AwFQ1T6GB9EF46DebNtEtMRoyKKxriPsue9Ez+ghcN+7
5+An3ZwlIXppRHGW/Fbe0rbbKsaCu8F1DqiBIvjL4FYNFh2DwitD7Ia5KB5D
Fqy2J34rCA6/cjoXYxtGd06cue7E53s7KTnByIXv0wmPQJH8HXsD03dRVBOy
ato/gKHpMWo5lAVh+bsTyAZirEYMJeYsjrPoYa3plU9EIAB9ZDfVIAU76xDQ
sp/7HgqM/nH7QyTpi9tzpRh9vsgZ7njvml+0rcSzmXhMvmBS+kGI9hMY/S+i
ZYJLznULNGIUNiZPoWYBS6l6ogGFGKPkTs84IFy7sS6hhviyoFBkk4j5gVBS
OfWi5mbRaZNPEhjBsGQ2rbvFkJDIiLdl/d7CHikyXgoLT0LT15bWM9xQfpJH
7YKbn0tiqR4QlJlkw6BcQ4KXVSX3L1j399+DmO5cc7SRbc8UxyBLEzXX1ngH
BCpsyMO2nTU8av+SFJ3qjacAwZFwpoadH9W7eM8F5Sv75F/yACdlehpi5cQE
U/ht4ykEQ5kyZqRFpr8dcMQKz8mrT8pMeBJC2hM5tLzmLJnvZgNDgh4xIJUW
YWix8hOLgUMVdOyVoNa/nYQ8C//W6TwnupbiuvLZht08DMboObEo+wVMuzuX
09I5WFhQJtPV1fV78gp2uCKHkW486Jp2gF/0QsJtRh5d7Mdv/bppbdelQVa+
O1ehXDxn7+wgEaX3abGB0f0CJlpfi2sJwla9gEYjKjGT7vO3O3VG4XD3BcD9
ZbryP6iPRXDiYKiN1peej1rCii3z7zsxFHkyun5E7pv87+SsOcbqjRpq4Ad6
RT9BYjpUIV8BqdL8c/VJQ24XWc79hPMcUBNL+2G+hRiDl0OYzs6KwsvInU6+
rRD5CRQcvlOfRgC6XIKMpoMR6vipy2qqhysAUdmjZWrj0oEh1yuBVQxAxld1
ay+tQROHyPZDKYMFOg33Iao+dD4JD9+ZIL/LGbI4Y4J0JvIuysotytziWWFI
4FTpPzBV5FMlEwklSeEXw0vgJ5LxGSYptu7Um+aTvblWTbT+wGyiBUjjCvHf
LeJrwzVeVwiChwjNp7bi+ugjq4H5yd9LhM3n2YdUG/wbJEyNj9KlIR5jkOdL
Xx0I7M7hSfBvXnOOpFDk5zP3y978693l5GiIl5exDZgAT9uNgCfSTvRqEPSL
tgl5sufmbpS6HOamgmV98EbX6aQ63uN7Z+/Ow2tkNNXwkWjUlRBP8gCiN+bD
LHbtH6p6jJswXXZj1D/952vM1dgifzPUmFe5/vZ58D3NSjgCKQpEHWC3XnAz
Y2xcatGhtlOziD8CzxqhkuS0ZA/GfZewt48TJZERDTy42ug/wZUScsz67OPP
Ynvm4JprCCvRxjwBcXXGGqBqNLkq6wLozVhNW2B51RH3UIv9zgQRs2EWRcVN
Vm4Nnv+H9FkG37s6XD8zJFj9LsiM+xUytnd8Vmm03Ar+k7GF0CpN2/n5+8X+
gWwC+NOQVmn/JfpHe3a7RfmZ+dOOhJ+1rODF7WWwVC9wg31o8IawfS/Tq+wy
ofXvw6QhXXeq0f70GX5vJQ/kZ2SzyTsXWNsbDZh2hziq2SrmounlqkpZwtoe
uzIMD5XVGFnDT6jkRWRSjuiujXliapusa9dWXJt7szazV17Zo/JQRrNx6Miz
nOBTtGnuj7h0MRXkVaugCR5mb9CZtV0y2n5jNPJp5f+4T2pEgdaetTGyhEIP
oSh0vLgWBXIfqwKOVUpRJVILPKLyn6xt9LcSiQIaCRk442ejWvy52osz7Ay8
6XfuwGEQFjVeIQaVVILbYYgp6y5UyBPHPjNqMiAhS9W4OQzAn5Qp6Bjz6Tfy
vTmaomrfH35IkgG6cC4oLp21qLsw5UbJhMNcQLpREJh8v/RycE+xgvjpve72
6XSP5IqV0MjNQf+IfS8+XsQ3NKtdY7cVUwg1NNTMODAfzDgzBB74ROYpVsMK
69VyVs8s1ILXQe8TVYRfYCDOGDjyIBzOvlFeV/cE0W9RNbWFG3tOimVJfznO
+uMteXA96EfG7gY9sFwkEDBTJ7f0two5pPSOvVgXF3rf0iZIlCJOkUyGdjSy
A4lF2epJrxAAGISJTx5Np41xOmYg1cUaiduIu5DZnMtxPwma6FHm66wJLz7w
QSbgapYosT5zXYC4a+3Y2/TpvfvLPYuVfAO5zFgSZQiw+vWyuflalYXlXY9a
s3Uh6/YfdpgKg4wmekJ6ZUXuHMdFzGXUahtiululay4EG2B6g94he1NvAv/0
48OdiBUMvH6AQsVeVYeAFP/DICd6i4wOI4md9KpBDcrV88r3Rd7b+os7DiUT
qFIds6z7ZEw0v1QA5a4EicOm1L/AAPYbl4L4ujJhVNffirzNIvZFIj+6db6l
nBpBpek0t5Wtk53C2iQ5AZxqQjzMXX1O/pMiuc8kllsC0C7rMfcRBUdd6fXj
zAhquTfIDGKUOh92x1mS4doVpjN9RkbkZ0a6uwzXCL1gCf2KZWxEsq/Lv5g+
U91yneVM/hCEnMycaS2k8jC7wsKAYa1JhT8Oifmiss99GfAxznB0XXdV6cL4
D1peZSOmszMjD3dd66QAxmosyoMvu7pA82hg0VLC9LFeetYtv5aNrHEeNQSb
sc+5SUVTVWlF5RuW0fQQNURf/JPhmdT3pAr5vdNjEh0y0JGTjzL2hxssSIi4
s2pK/8zRr7XAf+Q9qIq8GxWm7aw9aPSYvaYj1s9BL3OxHebDVFk624ix3Iu1
eBxMzx+uG3hbZGYwajlYZdYmLN02hlnqpPuTFyqF3XZ0QKn2Lt3dKM8RMnNW
/7h3DErGa8AF0dlQHqLl18s+fSYUGrmLIEVBbcW2FabjsCQ698ygx0+NFkqK
ga7lk0HIm2Xq2rYcc1WjpaJmejvBQhCTGtvkbMUfErNsd+3qJCV72texqb5T
gyoakRyHS0uQCLJApFeKg6jkWyaLZ/VDPAa7jhpH0lB8GkLxgDgrcIb/Thto
CXjgcTkYmY+AB7RIV1kubenL2cL+oacUHhcQRWkj+RpAA7sB1clgosR1/YGY
cYMAhgZF/fTPRyclGnjrK1pZTvnWshiigZdQEW4nlzGZFT4BjfEbDrLw3jlt
xNjUbUCDhnr8ehYGJLa+cDwF8176Bq5eoc22Nq6hO/Rswfotbsy89Nca8K9a
qrmd0QGofxibbVEbC8p88SUWf5AlGOJxJSV+TH3sgDN7ech73jGXxfwCE98s
uVu/2QDWhfCg7dIIbww8I7OEQRQCw0n+2Z0t8MRUmGwXrDhijSsvdRlO0ji9
7Ht7HxMLGyT/TZWqzszfbzTLuE5KoWE1/QRj6mGboVmB2KheTb5gIoXIDJBj
OioUfXo47O+sFU6IqY5Eu2Tsv/UU5kfMYEXWoJHavHZsbJ0F9YKPVz4SpIZC
SdTiXJ6UjViW/Nb31ux1n1nXeKXOez9jxPA3HllFO0wcmiR/U9FSxtxuB8y3
+ZY4zH6FuatK4pBZkGw/hI/qJ9FcKj+3yDKCWVJ1vs7m7b2qJ2iQ7lHfxYMf
WOywZrHomeN2COESJmzU6KBnu/gUgh2Mos574GJNcFWAGInZ5tbo953PxbQK
DPqo0Dk0qFSEfoTnW6puVD3x3f9rCM6P5I9DOELKYklLOwlPxJCOsrhRFKEO
naGeDd85nLa9z6P2cthr8rb73ZMGzZNhsvrt8InIzELttX9ltjXvK4KHN79p
c6wD+NEAiu+TzPrtqIBk1bMdOznQfcn6pkjTEdLRZqv4l75iNaTXpgk8MDZG
j4J6FMHziuOVkIyXAwnCtioMSrxXZg6CPdvddOfzrbPsqiGDHB9QoiIDly9m
8X1St3G704zZxxDiGAeeks+WFtg777l/v3eip4XMiooUoqI1y64JhtZWLnhf
RzAf6KPvgpPwOce5t06JLXFRCxaGMl21U3usBEqgnN24VSiHX+9fhyBjTnoI
DHxOYB/BvjJo6BTKNYQH3hSblYPpwmNtjGpIn8DK+XcIlD4kyjAMx27K7PYm
Wieyp8PHT3VeH0R9S0dhLrqk5WbxGflnaNDSD3TRYExyDOpg+xv6lV7k6UiU
iE99xfOScNLGLf2E22wmjCStEPLUtPJQQeHoCQDneUXgxSBBf+8Vi1O3NIhR
tbE74g14CSldIAysRhkYCE635J7t10ae+aYJCmoGqjR6KlEkDrmlXrrbWZd/
Xr04usoFJj1n9dyOmk0xQa7NRXBDrMtdmOYshq1Km1YTlV2pWSiBjFC9dbhL
KaDY3s5LSW9gMoj4dUjT3sMDheAfgio4Tf/H53p0KQiPXR/QXy+ZMOMj0el7
MF0vGK4bTO9XlKgy4wsZCZMTtz5Wrf9zrqnlcORhkheRcga9Qd90rKgGJFci
KJnW5gb1Cl3XC1eNvccDYFOsZQ2dPke8cE9xiYAv740XRViM4YCB7XQR8rcn
+5a6TiYVFv8n3xmJ2XkHfIV5HMaOVa+v28gygH/eq71gM+MSwoa3ZAxqBBTk
5xAv78sKnCuzgRzCjQ3xwKYKyffKIj7XkULrzyhVchfqYSdTK5J4V7EqpJKg
+ds3MkJllOs/AdUKLkYhT/wBhgwt4LtOG3bPxXfydASVf2k7ZjchbIa93bLX
sPCbNXUt8NZP49YnP+Qj7UWxlG4TWFexMRMgAInKxiMRy+SAQ6XkFITUA+qo
9jx/RkAjD+u9eQ8eIBmO7gQpl1W+r0NTJJnqp1aRDrhSpNRj7KJiUE3TntrP
pvAwzBGi1GyjJpgeMoQ1tOQAagB4ykghG4rJ2sEScsDZTWsDdUOflqmVqZ1v
NFVa3JuTVvf1ae0aihjzBJUD2ZG/rvO9udWTDr2b/usJxg5tA2d5XI1yDkW8
qM+mSG3r9054pSnxS3rkk31TT5d6bVTwxauBiTJq4703ZwiqQXNuOVuhamTe
HAeUjm8E6OtDCOupx0lb42Uy7fOVzDgzHH9nUoMY82KPNy6zmz1doPIyieI7
NCA5ds2IPNWquy7OfnJPa44N3zkIUFl5wr6CAMQWrGzx6+AoXD8k8aCbBaXE
+XVvF8gwOJxOry6kJZb5vI9riiRBSCo2ggsrC1nitK89sBuZZvjrZh8gb136
DQn6cRIHYqrMUZz0emrKzbCku/Vf+Pj/Vj+hVMhIalPqLPhNZEr37ZnZ8pP5
l7lQHeprWwUCcAWzsCLRBF7HgpLTNTOFTc2qF5LSLiMW4hAb8kNf5Sv9gEDm
ub9DCbWS4Ixv+cBFHhY+JFtgmkdXqmBjOkMsnxmpB4uJkPbSc8wpO41VGdcv
eifYxe4Bt/sGn1WYRqnHJdW1bRlUxgW5WJSrYAxFjNdJrKtWucnCx/2cGqXp
CfQT7Oi11h6ZhnBb8FPvMBDiSHVFmlW78dSrXU/hwNYTDdYXpqMbyUPrMhzb
L9yigWPXoD6XiBrknDlP46d0zWn5j7xoiKibQwcW/NWgtGtFDdl0UtMDRwyG
UTxLS+P9eoDAKmmOiF/ujdDPS/QLiVkKlK+DuXv41nghfRkwsr0DBeHO2Tj4
1+4clc8+FiGX7fIN69NkFfP/dh6qy6eWion84r7frfWyidG5BBvgAC38RlKu
NISCb8/ylcDLizMyMjOCqZnfrZu7BclrbgDZ0MSmtYg9BcXzXfRZTdDglKV3
T0SSwBDSsz2yrarBKypQMeSFuZZmUOYAnGwW978/FgLEqnwqFkVszansL3PY
5MhjfAdD7m2DAsBWd1Q21zYspL3Nm0niTgD5kiimx2YjxJmeUQZnZ2+bMI6N
vsLoc2I+1yeG2Kw3ti8iK1hSs5MKGPZA0zoVY4JV2GpG1zfRGtg39+3AuF4a
wokZxwqjT8rHFtslJZB3DSiN54rB4ggwImroePxgheWbx0nF0LqKUhxp7iqJ
dYi/Tc9RakA3zLQhkvK4XsM+Ir5/58u6KOLpdXpvDFgFbdP9KEOJ70eOYUeS
/nwNF8y0+MjLjl4m+uLdi7HDh/t4Bke5aew2/2HR5XBufWGJel+nsnEjmzMH
5DWBmsdBfXNj16O/tGAk3j0exEqSHKxCIIpjMiVmBT7pupEHUwRapwXyA0Dj
1uREbXOlM9Af6d+q1lv7p1Gcq3xoIHNaqSRAbqxk4ATekNpMazHXmx8fJEte
PnW+ibr5L8idWX2lYPSGeQ2Sv6zsk9ar34porZ7D5AfiaV+EAgxE6ZNdKSbk
AI0qhU6DEiZCzEpmh1qybPI65AGYPr69H40qsQNRxlLOns1bHgmaHDTATqYK
Ee17LEOIqUhzNs6g2ej/iFyi8RryGidEb4P7gZt8T13J94KhoJkavUqRjfaS
YezJBKi6FMGyyH36emMk+lwAtK2x1fKWDOHc0LQr4UaIZHp2+imkVSVL/iy4
nRuqBUryCsMOESUJyLgswHlpYe3t1WNePno0hZdIhELVH70AL8JqZ3hW/vrS
c9hpNAI25IDYGmXchmzWOBL6/Zzsx6bMiSG3/ljPN94jMEi7OOnNLm4F63xc
tnoA31gtIcHd8oscII5UNjxH6joCkM33cEpw4dKT7r2wl3aY1Ph5I6nDUpuP
rSzVyu+P6L1dDYnvFEHZRC/1qQ+3dzsSSvfDdS5wkHG3JyNp2KwEAoOBbcTw
6Q9Nrvt+ZoppjBqkJsM0oQc6+yG/WN5n4R5zXRGLI7Hf38ObcJzne7wM0hOO
Le2TE4m+pV6+9tGGJU3cSeYKCzRERuSuDBMigGjqaSxon7VCa6XYi0lCuzvq
423/6NMPN9XwUIvoAp1XKCbWoJjO85q0u9x5T0qWt1wytncRNW2hgk0tje6l
o57m3tgGvCqdYo3new+I8owhOQ8BRqZIYrQGzw0CxinxjTIsDp7x554TLrhA
cdcbYmIo7xBEPlCPSo8RyZ7u+a9xe2kJuFAVGGGE+Q2tlUxcuKWmIBvTJnB5
RAlKEVR1x+3RvQTXqzsezrV9z5qbG+BeQTzWmefMqtZQqLXujTrQ+fnY1syS
DJ7KjfUHwDxRjQf4DcoCKbd5s8MUlknTZK3SLAL7DqLI+dTv8lHRAH8zIhuM
AcQIDTXLMGR82oc4L1JbwGFUTcHg9mKfQWvYM4zOa+AYbMmqscD6PA/3qNN+
fuFSgEyYHsYStxssAL+CPrO4+OVGwdTaeh1qLPMmO2xDQwt0YH/k1xJ33jna
nVdS6VGaLjfy/jH23E9q6fnoR9QobDe0hsIXaBX8k5YaFK+u9bsIexW+ZkTD
IiM1JdQi90uVoDo9ekE4Yfqo1aWygXDsr3zFN2KCymiBYuI2x/PsI4k3M+Un
d0g3Rm6gaxmlAaD5cdxpjmNAcbn3zfxj3Q3IKwLbSrsx/BQBHXUJmwGdY9Lg
VYy2KfPjnavrlUIKGva+OH+CNJCEm9Y9+1z/KAzUGSX/Td48b9TRzi8/AKDK
DSxxgLetI5xUIyZ3BSjM0rdVbJMM6LGK43mfjejwqXy0jNaDr+O72lHD/pnc
iWbAAqwY2HlR6OF/z2rufvsPgovse18GE+8TBQlojmho0sbkO+PKxTzfIZAH
/mlPW7BsBlc4eP2mKy0XqOq02l359Se8cLUWMlFjjVmWwllWqmRy7noUi3ty
X36WDdNEr2RB2XL/kxW+428Lo6HGQrJ6VdiKyZoyVp6t93eLaNda8Aygjj7h
UhgRciWDlNq0ALYhzPev8K3m+RZj4sA2+J4JdPwv16gQ2fuk5rPdR1mGN1lu
sAN8xW+Iy/dcAcKO3BKB/i/+liEsWN+LLwNSuPQnBN+HRVw5eaUDe2aa8CTR
mlslag+ruX/ti8GF5/1m8KFQbb5+wQ0uVuQEyYwRm+lyyfLfpnh4436SNlaC
6cEaR1JavGratb5Vrri0Y8qosMOqG1sYTABn7GM0n8rXedJwM/aWWt6tZfnu
IJAYSo7sSqUxIECesPQz9lYeRKfDFLSUGFoGVuyqQY21+UtXuF8BPeLTfqpN
206gQqu+AyMlyejr2WFnBfCDmJj+RW2+19wYTxHkC+q8wQYAxI+BSnJ1/GTt
K9sQ8pZUI/ynBx6aThoTen2cPpDUn/wOGYfHaVlePp/wuXhDMCYCrgfCnFhm
RBUSRlDcR9399xh6YNesQ5fToDlGODXOQr554V3wXExM7ia++gmQWaycj0G0
F2bT53Wq0/1ExzwhrArYK5fzlFrbkwwDk9lE9C5irU18ZHVXlgWM4WrwUqN/
vhWJZ3q55PImwglNpzOg9U+dXx3OYq1m2BpH+giq95LH8nZwAj5WwhWHhRk2
Xg0t0OhljAR9nZ6ec4VMOfuMOGh6REhAMeP6T9SE7jicUkJ6Sigyqcm04+Y0
K05tb7xFv9Uj/HC6BXaCaVOQseHZDGABC5A/x/2LvGreYMf/hqEOsJ+hqH9o
TjQ4kQxF85v6zGaICkUk6ywvAXpbf36LefN723Mny3wvr2ztJxy3tvSwBp3N
g498PIKUqpQP9nVvb4QerzgPJDgCiATGJFGegx1aVsAKDNlGPVMXLZioV6EH
KkRGSmOOvDBH2/xjwTFDiHNUk/Z4IHSxE17AhVdszrNvoIcCJg7pqwm4ek7o
K5UvF9LWRCWvGlGZ8E4XTXbFNcdEwpyGKABccc6sQDKRkpu29IZeb9k+qemi
0zUWyOHGoF4733U09auqddRnDUv5t8r1AirtJxOsBb8R/CKIobIYaLlKjrkM
QiWdC7cd+D6KAw+x/cEfAfihF3ChZ9oA//feo4eooD+L1+n30OOAWmBWTMra
Use6VN6mnRy8iuFv+iJ42JrX+3cc0Nj29+UMn0nAOzi9dYGRSW+VpnL9k9/O
7MLSnW6sLybxsenHSyUXA5DoTXXaahPdf6X3QyQXTwRDF8E9E5P+HMyC76rM
ccf7V2bjqyUHtd+1sVINn65O+OsGUsmJQKrEEP1/4QDjmng0gl0Z2sf7pECa
9jxGJ+w+OamXXyj5et1J9mBObycvfk9hypKSM7rGVbazT0Az8B9rApeTIobn
dSC718kKY8X85T8ivH/81aTfODlCTeowy6lLeL57Yb3ejFWebqJX6ZvGvUnX
kteRjqCElUl7bZiHpUuPgrLN/Q7B/iBEB9uOnD5cjY4IfWqN2u2iT8GeRtOb
lj2Rpuduy0TO/0Th8eMVO2XJDkmtwpkAvYKmQ4cOL0vzrp3plWNJcg5mQ0Rj
uMI7QtwCUUFCqrlUyqqczPnrc/z0ESLC1Tu4TJGHoKenrLTZfIIv14rPEDX8
HSg4YPq50IGXbrKzBlhhqhlb7co8okaIHPEZIie54ovGNchCLjMojYqAL9i4
Iotc+2RtpWJM75HsHgjuXDuLsaMNnGW+WRDGtgIARy0LwP/ditT8K5qrXZc8
Z0BAQ7b4vI9cRsbz+8vFw4fsF3ElIYB9bZKOUvTJMVeG0E+BOnT2anAH28j1
YxwGrer+NPRWxtq52dWvgplR93RTbdG8xjWyS6052lPiNqA+KlmRY+4ETrBj
K+0LZ+EUFBmIf+HKQchOvWEaSgK7W4SEUTCyxPiS00gAepPiJEJ1lXOHzjTm
r5VlwB9QFQDtnoFHT9aZrhcPrAqi4dglw1uopbfU24f9tQx8uBemIvo/irNC
786keS32HCv8O5d07Pbr26NaE+0JY5aXdX8Ks2r8zlFvVvrI52iENB8Mc9or
Tm+0TDgvWjSR8PeODrz9qbNjpkoLjtIjL8L7xZERWeppm9UzQlFfGukDNMdZ
DRC6gFMMY0BNg7zsG6lTbAZ+SPcNeOzlmb7dR7+QdNQd/68OI9Z4SDVIh0sa
U+ogHqh/B5ZXywqcCpMYvANIrM/yJI395DDzeim2gPt+hhitKAjwHiY8N6TV
gEi8BOKXq14UaDUwD/BEpEIa84TmD7uqtan9Vjj3frvtUAdUB/MRIZ00JOdh
3pHu5wEyqiql3z7IawG/MeO6VaxefFsXvkSzETRqPiFFJf29pMGxjHb8w0y0
Lq+eONZUtULAEvJhDxKNX7YfO4KjVDvLFqS/3ctYunwMonJjtPZOueV49ObK
Jmtk0aTj6Oc4YJuZ04qSkfMQSgmFzKQ1xSGXVNUW4DtDmyG4pyr85zlVG2j/
OjXslkDS8aUWP10Mm0n1MxKIpY4UV0DaficioL33K+y/PhmCKLbrIL5tMc/t
3ajoj+6mkQGENCW5OMxfI7XP2Y0Sa4vEbKB96444L73BvwA7LMeAcoDFwpT/
LDJ1zioKFpdLhNbkmPA2dsvQOHgDfVamqb+vOLRjF1JbhQieYZHhhaBi2BN3
JkFWisKasYfHOvkGF5A3RVraQx8y+ScOqqcSiPvYwYLuEfaqs3rGVW7UDfsx
zCQg11EqJtY1i7RCIeiuV8U04G2GMFidXVnPZuVlqs+dRzdkPlaXDCFpznc6
ImzB2zKDMTiqgnj0hQ98Gjxk1K60G5+scdfQnZpYf63yCC6AvJf1tQUx0h/g
wcth3DSBSiUPEzucIYvqqhcj7HCxHY9TLwyjOT6o5OXH8zSbU5lXm5vASV6Z
WT5+q6Rct+MlqjBrm4mmJToS/jbZSd0uPMJJ2CTogFwaGvy+1CLVTfH2rHCD
pFQKT7Xl52Rxmd0Lcnj1I/zsc17xfqGcUygl8S09Cyzy6ziyJJAtg3xFMYvB
3oFDmYykIIYxzJCQkYof5C1KopaKcsKzxT7vqp0vTGgE8d4Cyz1f4N21kdK3
dwj8N2VSrDUlGaRNSoJH1RGjrYBM4+5GlODFlYeOo1SZ48jPbFBBGp+EK4xP
q+cOx1cpNF9nxdggfjRalpQWnbnEwgkEKDq3RrCiHgmfB10U8mP1MhTjJLMq
uhnhKJkbl9pueb6fJ6h650er/g5/XtDmi6218rr03sYrEBIWQ7O9pnfZTAij
OlbVEVd8mfxSH0zHC1YPxuDosrAmxay3tC3zaRLvCABqaltW3hkL7toXTRW5
Y/pW2kvTfWNYSKkyhmV47//DGV5jEgFVjoOrFNFcbHGDfItQ2QnB8gt/LWNB
7f7/yCVTm9A5PGU3my+oyWOq8rUf1UFvBS6cV04OuOByTvWgZeCY7/+AsWg0
gcrcw+2n5fj11LxryxeNG+40/wyw1/KYnP8l8ZSaTb7qHj5zbu2f7DDbWG8E
zcK2oFdiwFusKUxrWe8QoRgjekq2hAX2nw0HtKDbBxePqL23fmED3qMcBeID
pECNvGO5mcZnu4SEKYn6QKV5RVBpiu7cYjArYe60k/VHivfjdKdPH6KLaMKr
CgnTFF8GiK+erRN3QGH8B2YVgQZD0sutKkWp7UEdhZBqvi9pPo1h7qw2mqXm
Nyqo7XI08W/Fd4kZVEY8c0MPk/I7GqPhGOtP9JQFBmKwhWigsPZQZwbyS6vU
Hiz/0HcZD4ZSIkilwJ7/q6O/9r7D2OxlZZBtWCCjjVa56Nkwrqb/Y7cHgMMq
ghxsQ82tlmj+mkmeSWsEkjmu6qJ2mEoZvFR/ySsOGgCTq+0WiJMz9ZlhQu7y
dawnW9NJbXYmgvVDJYpPzD+4nPNyZrURWNPxzr98KEnSrDUENpmBvcnKS+Sg
Cc+PFXLFetLBsTPIozUmmdlkx9h01ZK8MirhvuFltbpvJGVXdoegpWcyGeEg
aYtnV5qxNLOj2L6pHCF3ufNSMaZfoEsjO9vrWDTt41OXkS98I8H2cTvCuzJd
tqNH5n05iaSCzdvtanQM4jL+1zmM7iACkf+EqnX1qxuNBX5H3qW/SMenGDgO
xYXXfraaOUAkVhu00IBJGnGZNHk/3SvGnPlgwNersqS2fA6b40VNUO1VQ1oJ
nG5Nyj9IOdI6KedoZ5aDNWid8FlZNqxcoYJWS9iKd9yql2ig05n18jZZt1Xb
3zX5TXCK4ZqaRMq3Sp7KHkJhE78cJJ0mITQ2iPdqOE8HsD0P+qlu665GgQTu
KMHZgU/6/nYQk2pxGmAdZavyLXGvDsNhZQKbNo2ZVsm4iFPs7UO9tSKaaia6
/0OrRqSl9do9LaGWP+ORqIWArZaEfBFfd5p8cIdQaVd4TrUIoCHIDmSHPOG6
XzX3upxyu26xz+f9YrRyjdtx/7SL8ajS2Ptjcs0H2xT1uFVDKcZq0OMumpG2
pQY6M7i0WVfp8aVFoxRyhMjlbDelafuwu7a7H79mXyWuif0KFTEokOIksYR/
JyvO+8Zo9G/ytzwDmHVNH98KHaT4QcHnYSzU8oBI0BEJBavIEd1fYcnEFX49
RwCpKQDYMWC4A5nXJ0WGrSmkOEcoXaZAh//7Gn0HP5aCDPr0uBCK8DFP2hXm
5xUozf2+ED1ulncVOE3A8cOT4D0MQev20zGQvlx3gUbZsX71wHo/90VEehTP
aHNvzFPL7VZwnd1jLD2I2G99JwkxfLckBSOHa3Ug2V963xSp8B+ko9yFo2jN
Jjf/ZQmCmySgM3parlGxlHMr/RHee55/ohxVPd/3qxaA7CuYAfy4eefG+uAh
NZmYonx7LgaP9vLCsXmfO53a3JLm/qLmGya/gDYz/CnPgZcf3bKJBhx+ZqPq
6AkQuPVxrocIJBcDU082eoTPwonROKvxOHPBwykm1GeOH4rE7hSlqOORfYad
ONJgx31sJictcT/mb3Hz2CyX9dF0zMReyN/w2vGpkq/zoBn+h075gueCsa+o
N+Kz0JcpQkYq8qNwHlGM7VJ8R/i3QilGZZ1uv781D8RRAYPecm9fr7xUMTe2
JxAmHJDiQMF4BcEc/rY7+/m7xL/aHtpZVk/J3ZoOfeP/EmFAgqmsl4hXhQiq
fax00tjahqcJ2h9bvvyBDNLGEM9UUPUrYwOKY+PcXsQTU4QBLOCKCoGT61Bh
AAUgp4HbilybvLrk4M5mT/zy/SKs7Wq4fT/HtPEkfHPT+u9C26JnDnYSDFqY
uZIncwF28/YprhSXgLrX3Tv5zm/XHu7NWe+pWMLof9rweSrdI1lbjApvDhIJ
h0SpyTpRvHI2EHGLMs1uDjL9TUUiWfwUyAHTO7gdBNXyvaymE9gY2+vY5WPW
U2hAOwsrfbODyfi+/3k4dFKpryFpmobnv5o79y2Ef5wF0g0igxIwMv0eRaU1
Nf7NUTjH58spsiG4AU1O9xQfUXWh26LnxtopOJg5T5CZ1YYrHsBcSSgxoVdA
j/FUls2XBVNWCVgTMFCbcvxbCgkTQHFX1CUMfudE6rwOa0bQ2acVU2Oin+r8
88NJABY6f3HcQI5XSrp8Wn8XC+02pRymuD94WoQQMGW8F+uQcSwCaQDNKJvI
1etsRnXS30VuAMpPsTTagAkdJ8MdT5gXu2D8V19ROqjAHzDURLKjI/8For0M
MTTOdsyTajzX0kP/XzsRBfNNHiiDqJv5Rls+m/wJ1My4/MSvpF+pJL2LZPu/
7hDfxEXi8KoRdNop4U8lNiP/PSbTfeQZNx864ygPTEuftPl9kj/MdP/MkPDe
6k+RNUMUw+KmsR9Bv1PHdDkxug6YGXN12MEAb7+i4U4ONA5r+OwU78yuyPjM
pTzV16ZtjxpijPAtu84ddTA5/3+/QJyK+SQULrjkibIoQeRVQ5bI6KeOSNav
tsnRGOkWY3o/DRwUI2313MT3P/+8G4EH4AWAqKluQBVNqAt144giUJezrIhN
nq6Q3MsVFV/xQWU/T23vG/LUmvoITekYP23A7WG6JKjlzmZORFKXQuOH9cNv
8EYnoSlSrJhkgIfxyAmjRxb3HqYoa4fZg2OcsgrBw2OUBk/6iLE3EVvCWQ47
qZb6jiQ+In9QJxtt1Bs9vspO5C6CUlwlKX3vhFyAEBTSiHKTTJzIX5GovAvb
dlil5fDVRgdf/QqYYdNaJxy5qkgKHcDoLw7E5DFGV48vrXUy2YlDVPnHASHO
tLvoMkyhhEp/5BusgbXWoMIC34tz4TH+cJAOOnGcvCCebZJNhJICi0m02mt8
6jftvBS7+1n+jaDs3U1NqfaA8f9N+VycW5CwOsSbAg2eHCO0oIzrIr3eG3nn
RvCHxR8qaif0ED3JvxTT7P7GHxnfuJEU0a7MycnaqWJJI3HacMJYQHhy0QT3
NIk8RIcMIgknyosYdVDi+F1iWpZjmPeYedIlNlG4ZgWGTaT9XTrFlcoQrylz
wD7aGPnXSs0TGXwnNcoXtOvXZkfOtYVcho2ad45LNN26hSxHYq/7Nu9xB4h6
LLzGiyBlxYfMt4pErmqo90pXc29NZTOsgffPTEbosxC9tCZQBofy1+I2gjdP
iLesnW/rrlidKrLg61TGo1qC2hDM0X7+jDvNJVGazSlK7XhxMMZV8qGxt/e6
yU0dJzPy4Uz77p51p1HPIiCjFfrfU93JEvuTjOqK43hahprQDoWIO8knC9Ce
scvVl+S8wkIVi9lH1jT81a41HOk/PU/EPCfOCpCjG62zgic8INrDk+CbXAVL
ilWSxKnR7S9rROthl9dwso5NgD6vLDS7pCgkFWhTdnNROqI7cVbNIz5Flews
QQgvTJ8rFVzFF1iNSss/GpblzcLBJd9INF0ddcAyQ3lJjpTswNSlorqohV75
zClUOsH+ypaoH7Q7fJ5+5q2SPhBpi232KpepTl0WPolzblAWahA5gZGI2P8+
Ht1J7XQwylQnARaw/hHhsUlQoZg7xn/Tf7UX2bwT4PEsr8b/1II1P5sLP/YC
okvAFbyVgsbXg6Lw2tFfRnqvuzGx4M5I7xIiYpIZOIDBgjklWBTdcLhnRCXN
aSx23smzIWkXMDF8OtKFxfD45pcJYB9lf/mOlhNj7BTGAGgHhPXZAEBTXUaD
9c3iDYzM/PfcDYISlQjNicMeqYtZM4RfoaLl7zvU8bjSlVww8exKEM/3y8aE
W8DZYympXLq6FPEMWINei13myBTXU1JuHmtpFbkxXNkHoui8gcSiWnfS4i5m
TC1qv86NT+02YzEF

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "OJXsOzX3SCOyhcBXS9yryN9cWQxQkhDHUr4mzQikLKNKnB6JkSYY9xNnmYkvVOJ5f3SnsxLM71tWjwpqmyTCVkTt4jikDmXDCnl6lQn2TVy78ivgbebFE/F7GUr3Z8AASPmtz4v12cD/Cz7nTJMTG81IGzEoV1S4KsV3MBcbB+1TqTshtjzQ4oMMPpNw9ltjOjjqx8CktvtqLiQWjnKfQh8i3R/5yQlzObBDq+VCqANlykTDX90l/EChOZyM2vP2LPtHKdTejov5NWYnpITxaU4mVC0qHRZWMw311CSPr2DthD+mQpU6WB0IW0Q/RSRVGukl/zoGSJK4WPzZBsbx0qQYZKoOugYWEzdhvyM9sRbw8X8It1PqMRIkjL2HSiU2Yamr9tujeh3nZc8bAS2APHiTCghwu1UxljKiPz93UDwPV04N10QIv52NKTBZZFxBZEcn16ksA0USMMfkVi56IRF3SVObWZkPdB+eTvGsXvilaS9Z+DoKm7ewTiLUp4m2ltYuN3vHs/IS7T00K8KNnQzXnqfgjutEQ1sUj6JHTqjHml3CSrEe1oCyfTnGdhX6w8N4YMxU7nS157ZrwgAOiQc1YAFZZMAljXxwHvd5kOTJAOxcok27gjNW6qiHriXmrIpdaJtyjanuDAv4dN65QI5NWp+t3GDSAifEFcfwfhGXd3y4ZQwffvJLAAyKcdTlQgfJqXgaeK27hhml4j+dtoKIeF82AkAZFUOZQEG7rzb4w/nX6GHDXSIFO4jK3VlGo2LftMj45bOOKgfCDFAgtBU1L2P36etR5cT9dZ5PSpLxdOOdTIWtgi9kZ1NbD33gDcr0hq2g1R5UMiIhFQLyoKkbGvIiZPAfTzySQH65nPorjqLPwAgNawFc3UnRn7ch8dPTUo/KBPppziAa1Nx/gRJhFwsNYd2EJkSQr40IHJcV4cTS9rdxboidvaIUo4Bf6F2bsV9YjWFrHgx0LhtFnBSyWuSD9wxmkIEqTEDuB5RJtaqjrDhuZnZ3Z3mxFqAT"
`endif