// address_decoder_top.v

// Generated using ACDS version 23.4 79

`timescale 1 ps / 1 ps
module address_decoder_top (
		input  wire        csr_clk_clk,                             //                     csr_clk.clk
		input  wire        csr_clk_reset_reset_n,                   //               csr_clk_reset.reset_n
		input  wire        mac_clk_clk,                             //                     mac_clk.clk
		input  wire        mac_clk_reset_reset_n,                   //               mac_clk_reset.reset_n
		input  wire [25:0] slave_address,                           //                       slave.address
		output wire        slave_waitrequest,                       //                            .waitrequest
		input  wire        slave_read,                              //                            .read
		output wire [31:0] slave_readdata,                          //                            .readdata
		output wire        slave_readdatavalid,                     //                            .readdatavalid
		input  wire        slave_write,                             //                            .write
		input  wire [31:0] slave_writedata,                         //                            .writedata
		output wire [19:0] multi_channel_address,                   //               multi_channel.address
		output wire        multi_channel_write,                     //                            .write
		output wire        multi_channel_read,                      //                            .read
		input  wire [31:0] multi_channel_readdata,                  //                            .readdata
		output wire [31:0] multi_channel_writedata,                 //                            .writedata
		input  wire        multi_channel_waitrequest,               //                            .waitrequest
		output wire [13:0] traffic_controller_ch_0_1_address,       //   traffic_controller_ch_0_1.address
		output wire        traffic_controller_ch_0_1_write,         //                            .write
		output wire        traffic_controller_ch_0_1_read,          //                            .read
		input  wire [31:0] traffic_controller_ch_0_1_readdata,      //                            .readdata
		output wire [31:0] traffic_controller_ch_0_1_writedata,     //                            .writedata
		input  wire        traffic_controller_ch_0_1_waitrequest,   //                            .waitrequest
		output wire [13:0] traffic_controller_ch_10_11_address,     // traffic_controller_ch_10_11.address
		output wire        traffic_controller_ch_10_11_write,       //                            .write
		output wire        traffic_controller_ch_10_11_read,        //                            .read
		input  wire [31:0] traffic_controller_ch_10_11_readdata,    //                            .readdata
		output wire [31:0] traffic_controller_ch_10_11_writedata,   //                            .writedata
		input  wire        traffic_controller_ch_10_11_waitrequest, //                            .waitrequest
		output wire [13:0] traffic_controller_ch_2_3_address,       //   traffic_controller_ch_2_3.address
		output wire        traffic_controller_ch_2_3_write,         //                            .write
		output wire        traffic_controller_ch_2_3_read,          //                            .read
		input  wire [31:0] traffic_controller_ch_2_3_readdata,      //                            .readdata
		output wire [31:0] traffic_controller_ch_2_3_writedata,     //                            .writedata
		input  wire        traffic_controller_ch_2_3_waitrequest,   //                            .waitrequest
		output wire [13:0] traffic_controller_ch_4_5_address,       //   traffic_controller_ch_4_5.address
		output wire        traffic_controller_ch_4_5_write,         //                            .write
		output wire        traffic_controller_ch_4_5_read,          //                            .read
		input  wire [31:0] traffic_controller_ch_4_5_readdata,      //                            .readdata
		output wire [31:0] traffic_controller_ch_4_5_writedata,     //                            .writedata
		input  wire        traffic_controller_ch_4_5_waitrequest,   //                            .waitrequest
		output wire [13:0] traffic_controller_ch_6_7_address,       //   traffic_controller_ch_6_7.address
		output wire        traffic_controller_ch_6_7_write,         //                            .write
		output wire        traffic_controller_ch_6_7_read,          //                            .read
		input  wire [31:0] traffic_controller_ch_6_7_readdata,      //                            .readdata
		output wire [31:0] traffic_controller_ch_6_7_writedata,     //                            .writedata
		input  wire        traffic_controller_ch_6_7_waitrequest,   //                            .waitrequest
		output wire [13:0] traffic_controller_ch_8_9_address,       //   traffic_controller_ch_8_9.address
		output wire        traffic_controller_ch_8_9_write,         //                            .write
		output wire        traffic_controller_ch_8_9_read,          //                            .read
		input  wire [31:0] traffic_controller_ch_8_9_readdata,      //                            .readdata
		output wire [31:0] traffic_controller_ch_8_9_writedata,     //                            .writedata
		input  wire        traffic_controller_ch_8_9_waitrequest    //                            .waitrequest
	);

	wire         csr_clk_clk_clk;                                                                      // csr_clk:clk_out -> [master:clk, mm_clock_crossing_bridge:s0_clk, mm_interconnect_0:csr_clk_clk_clk, multi_channel:clk, rst_controller:clk]
	wire         mac_clk_clk_clk;                                                                      // mac_clk:clk_out -> [mm_clock_crossing_bridge:m0_clk, mm_interconnect_1:mac_clk_clk_clk, rst_controller_001:clk, traffic_controller_ch_0_1:clk, traffic_controller_ch_10_11:clk, traffic_controller_ch_2_3:clk, traffic_controller_ch_4_5:clk, traffic_controller_ch_6_7:clk, traffic_controller_ch_8_9:clk]
	wire         master_avalon_universal_master_0_waitrequest;                                         // mm_interconnect_0:master_avalon_universal_master_0_waitrequest -> master:uav_waitrequest
	wire  [31:0] master_avalon_universal_master_0_readdata;                                            // mm_interconnect_0:master_avalon_universal_master_0_readdata -> master:uav_readdata
	wire         master_avalon_universal_master_0_debugaccess;                                         // master:uav_debugaccess -> mm_interconnect_0:master_avalon_universal_master_0_debugaccess
	wire  [31:0] master_avalon_universal_master_0_address;                                             // master:uav_address -> mm_interconnect_0:master_avalon_universal_master_0_address
	wire         master_avalon_universal_master_0_read;                                                // master:uav_read -> mm_interconnect_0:master_avalon_universal_master_0_read
	wire   [3:0] master_avalon_universal_master_0_byteenable;                                          // master:uav_byteenable -> mm_interconnect_0:master_avalon_universal_master_0_byteenable
	wire         master_avalon_universal_master_0_readdatavalid;                                       // mm_interconnect_0:master_avalon_universal_master_0_readdatavalid -> master:uav_readdatavalid
	wire         master_avalon_universal_master_0_lock;                                                // master:uav_lock -> mm_interconnect_0:master_avalon_universal_master_0_lock
	wire         master_avalon_universal_master_0_write;                                               // master:uav_write -> mm_interconnect_0:master_avalon_universal_master_0_write
	wire  [31:0] master_avalon_universal_master_0_writedata;                                           // master:uav_writedata -> mm_interconnect_0:master_avalon_universal_master_0_writedata
	wire   [2:0] master_avalon_universal_master_0_burstcount;                                          // master:uav_burstcount -> mm_interconnect_0:master_avalon_universal_master_0_burstcount
	wire  [31:0] mm_interconnect_0_multi_channel_avalon_universal_slave_0_readdata;                    // multi_channel:uav_readdata -> mm_interconnect_0:multi_channel_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_multi_channel_avalon_universal_slave_0_waitrequest;                 // multi_channel:uav_waitrequest -> mm_interconnect_0:multi_channel_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_multi_channel_avalon_universal_slave_0_debugaccess;                 // mm_interconnect_0:multi_channel_avalon_universal_slave_0_debugaccess -> multi_channel:uav_debugaccess
	wire  [19:0] mm_interconnect_0_multi_channel_avalon_universal_slave_0_address;                     // mm_interconnect_0:multi_channel_avalon_universal_slave_0_address -> multi_channel:uav_address
	wire         mm_interconnect_0_multi_channel_avalon_universal_slave_0_read;                        // mm_interconnect_0:multi_channel_avalon_universal_slave_0_read -> multi_channel:uav_read
	wire   [3:0] mm_interconnect_0_multi_channel_avalon_universal_slave_0_byteenable;                  // mm_interconnect_0:multi_channel_avalon_universal_slave_0_byteenable -> multi_channel:uav_byteenable
	wire         mm_interconnect_0_multi_channel_avalon_universal_slave_0_readdatavalid;               // multi_channel:uav_readdatavalid -> mm_interconnect_0:multi_channel_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_multi_channel_avalon_universal_slave_0_lock;                        // mm_interconnect_0:multi_channel_avalon_universal_slave_0_lock -> multi_channel:uav_lock
	wire         mm_interconnect_0_multi_channel_avalon_universal_slave_0_write;                       // mm_interconnect_0:multi_channel_avalon_universal_slave_0_write -> multi_channel:uav_write
	wire  [31:0] mm_interconnect_0_multi_channel_avalon_universal_slave_0_writedata;                   // mm_interconnect_0:multi_channel_avalon_universal_slave_0_writedata -> multi_channel:uav_writedata
	wire   [2:0] mm_interconnect_0_multi_channel_avalon_universal_slave_0_burstcount;                  // mm_interconnect_0:multi_channel_avalon_universal_slave_0_burstcount -> multi_channel:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata;                               // mm_clock_crossing_bridge:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest;                            // mm_clock_crossing_bridge:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_s0_waitrequest
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess;                            // mm_interconnect_0:mm_clock_crossing_bridge_s0_debugaccess -> mm_clock_crossing_bridge:s0_debugaccess
	wire  [16:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_address;                                // mm_interconnect_0:mm_clock_crossing_bridge_s0_address -> mm_clock_crossing_bridge:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_read;                                   // mm_interconnect_0:mm_clock_crossing_bridge_s0_read -> mm_clock_crossing_bridge:s0_read
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable;                             // mm_interconnect_0:mm_clock_crossing_bridge_s0_byteenable -> mm_clock_crossing_bridge:s0_byteenable
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid;                          // mm_clock_crossing_bridge:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdatavalid
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_write;                                  // mm_interconnect_0:mm_clock_crossing_bridge_s0_write -> mm_clock_crossing_bridge:s0_write
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata;                              // mm_interconnect_0:mm_clock_crossing_bridge_s0_writedata -> mm_clock_crossing_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount;                             // mm_interconnect_0:mm_clock_crossing_bridge_s0_burstcount -> mm_clock_crossing_bridge:s0_burstcount
	wire         mm_clock_crossing_bridge_m0_waitrequest;                                              // mm_interconnect_1:mm_clock_crossing_bridge_m0_waitrequest -> mm_clock_crossing_bridge:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_m0_readdata;                                                 // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdata -> mm_clock_crossing_bridge:m0_readdata
	wire         mm_clock_crossing_bridge_m0_debugaccess;                                              // mm_clock_crossing_bridge:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_m0_debugaccess
	wire  [16:0] mm_clock_crossing_bridge_m0_address;                                                  // mm_clock_crossing_bridge:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_m0_address
	wire         mm_clock_crossing_bridge_m0_read;                                                     // mm_clock_crossing_bridge:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_m0_read
	wire   [3:0] mm_clock_crossing_bridge_m0_byteenable;                                               // mm_clock_crossing_bridge:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_m0_byteenable
	wire         mm_clock_crossing_bridge_m0_readdatavalid;                                            // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdatavalid -> mm_clock_crossing_bridge:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_m0_writedata;                                                // mm_clock_crossing_bridge:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_m0_writedata
	wire         mm_clock_crossing_bridge_m0_write;                                                    // mm_clock_crossing_bridge:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_m0_write
	wire   [0:0] mm_clock_crossing_bridge_m0_burstcount;                                               // mm_clock_crossing_bridge:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_m0_burstcount
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_readdata;        // traffic_controller_ch_0_1:uav_readdata -> mm_interconnect_1:traffic_controller_ch_0_1_avalon_universal_slave_0_readdata
	wire         mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_waitrequest;     // traffic_controller_ch_0_1:uav_waitrequest -> mm_interconnect_1:traffic_controller_ch_0_1_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_debugaccess;     // mm_interconnect_1:traffic_controller_ch_0_1_avalon_universal_slave_0_debugaccess -> traffic_controller_ch_0_1:uav_debugaccess
	wire  [13:0] mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_address;         // mm_interconnect_1:traffic_controller_ch_0_1_avalon_universal_slave_0_address -> traffic_controller_ch_0_1:uav_address
	wire         mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_read;            // mm_interconnect_1:traffic_controller_ch_0_1_avalon_universal_slave_0_read -> traffic_controller_ch_0_1:uav_read
	wire   [3:0] mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_byteenable;      // mm_interconnect_1:traffic_controller_ch_0_1_avalon_universal_slave_0_byteenable -> traffic_controller_ch_0_1:uav_byteenable
	wire         mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_readdatavalid;   // traffic_controller_ch_0_1:uav_readdatavalid -> mm_interconnect_1:traffic_controller_ch_0_1_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_lock;            // mm_interconnect_1:traffic_controller_ch_0_1_avalon_universal_slave_0_lock -> traffic_controller_ch_0_1:uav_lock
	wire         mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_write;           // mm_interconnect_1:traffic_controller_ch_0_1_avalon_universal_slave_0_write -> traffic_controller_ch_0_1:uav_write
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_writedata;       // mm_interconnect_1:traffic_controller_ch_0_1_avalon_universal_slave_0_writedata -> traffic_controller_ch_0_1:uav_writedata
	wire   [2:0] mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_burstcount;      // mm_interconnect_1:traffic_controller_ch_0_1_avalon_universal_slave_0_burstcount -> traffic_controller_ch_0_1:uav_burstcount
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_readdata;        // traffic_controller_ch_2_3:uav_readdata -> mm_interconnect_1:traffic_controller_ch_2_3_avalon_universal_slave_0_readdata
	wire         mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_waitrequest;     // traffic_controller_ch_2_3:uav_waitrequest -> mm_interconnect_1:traffic_controller_ch_2_3_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_debugaccess;     // mm_interconnect_1:traffic_controller_ch_2_3_avalon_universal_slave_0_debugaccess -> traffic_controller_ch_2_3:uav_debugaccess
	wire  [13:0] mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_address;         // mm_interconnect_1:traffic_controller_ch_2_3_avalon_universal_slave_0_address -> traffic_controller_ch_2_3:uav_address
	wire         mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_read;            // mm_interconnect_1:traffic_controller_ch_2_3_avalon_universal_slave_0_read -> traffic_controller_ch_2_3:uav_read
	wire   [3:0] mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_byteenable;      // mm_interconnect_1:traffic_controller_ch_2_3_avalon_universal_slave_0_byteenable -> traffic_controller_ch_2_3:uav_byteenable
	wire         mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_readdatavalid;   // traffic_controller_ch_2_3:uav_readdatavalid -> mm_interconnect_1:traffic_controller_ch_2_3_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_lock;            // mm_interconnect_1:traffic_controller_ch_2_3_avalon_universal_slave_0_lock -> traffic_controller_ch_2_3:uav_lock
	wire         mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_write;           // mm_interconnect_1:traffic_controller_ch_2_3_avalon_universal_slave_0_write -> traffic_controller_ch_2_3:uav_write
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_writedata;       // mm_interconnect_1:traffic_controller_ch_2_3_avalon_universal_slave_0_writedata -> traffic_controller_ch_2_3:uav_writedata
	wire   [2:0] mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_burstcount;      // mm_interconnect_1:traffic_controller_ch_2_3_avalon_universal_slave_0_burstcount -> traffic_controller_ch_2_3:uav_burstcount
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_readdata;        // traffic_controller_ch_4_5:uav_readdata -> mm_interconnect_1:traffic_controller_ch_4_5_avalon_universal_slave_0_readdata
	wire         mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_waitrequest;     // traffic_controller_ch_4_5:uav_waitrequest -> mm_interconnect_1:traffic_controller_ch_4_5_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_debugaccess;     // mm_interconnect_1:traffic_controller_ch_4_5_avalon_universal_slave_0_debugaccess -> traffic_controller_ch_4_5:uav_debugaccess
	wire  [13:0] mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_address;         // mm_interconnect_1:traffic_controller_ch_4_5_avalon_universal_slave_0_address -> traffic_controller_ch_4_5:uav_address
	wire         mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_read;            // mm_interconnect_1:traffic_controller_ch_4_5_avalon_universal_slave_0_read -> traffic_controller_ch_4_5:uav_read
	wire   [3:0] mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_byteenable;      // mm_interconnect_1:traffic_controller_ch_4_5_avalon_universal_slave_0_byteenable -> traffic_controller_ch_4_5:uav_byteenable
	wire         mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_readdatavalid;   // traffic_controller_ch_4_5:uav_readdatavalid -> mm_interconnect_1:traffic_controller_ch_4_5_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_lock;            // mm_interconnect_1:traffic_controller_ch_4_5_avalon_universal_slave_0_lock -> traffic_controller_ch_4_5:uav_lock
	wire         mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_write;           // mm_interconnect_1:traffic_controller_ch_4_5_avalon_universal_slave_0_write -> traffic_controller_ch_4_5:uav_write
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_writedata;       // mm_interconnect_1:traffic_controller_ch_4_5_avalon_universal_slave_0_writedata -> traffic_controller_ch_4_5:uav_writedata
	wire   [2:0] mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_burstcount;      // mm_interconnect_1:traffic_controller_ch_4_5_avalon_universal_slave_0_burstcount -> traffic_controller_ch_4_5:uav_burstcount
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_readdata;        // traffic_controller_ch_6_7:uav_readdata -> mm_interconnect_1:traffic_controller_ch_6_7_avalon_universal_slave_0_readdata
	wire         mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_waitrequest;     // traffic_controller_ch_6_7:uav_waitrequest -> mm_interconnect_1:traffic_controller_ch_6_7_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_debugaccess;     // mm_interconnect_1:traffic_controller_ch_6_7_avalon_universal_slave_0_debugaccess -> traffic_controller_ch_6_7:uav_debugaccess
	wire  [13:0] mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_address;         // mm_interconnect_1:traffic_controller_ch_6_7_avalon_universal_slave_0_address -> traffic_controller_ch_6_7:uav_address
	wire         mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_read;            // mm_interconnect_1:traffic_controller_ch_6_7_avalon_universal_slave_0_read -> traffic_controller_ch_6_7:uav_read
	wire   [3:0] mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_byteenable;      // mm_interconnect_1:traffic_controller_ch_6_7_avalon_universal_slave_0_byteenable -> traffic_controller_ch_6_7:uav_byteenable
	wire         mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_readdatavalid;   // traffic_controller_ch_6_7:uav_readdatavalid -> mm_interconnect_1:traffic_controller_ch_6_7_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_lock;            // mm_interconnect_1:traffic_controller_ch_6_7_avalon_universal_slave_0_lock -> traffic_controller_ch_6_7:uav_lock
	wire         mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_write;           // mm_interconnect_1:traffic_controller_ch_6_7_avalon_universal_slave_0_write -> traffic_controller_ch_6_7:uav_write
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_writedata;       // mm_interconnect_1:traffic_controller_ch_6_7_avalon_universal_slave_0_writedata -> traffic_controller_ch_6_7:uav_writedata
	wire   [2:0] mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_burstcount;      // mm_interconnect_1:traffic_controller_ch_6_7_avalon_universal_slave_0_burstcount -> traffic_controller_ch_6_7:uav_burstcount
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_readdata;        // traffic_controller_ch_8_9:uav_readdata -> mm_interconnect_1:traffic_controller_ch_8_9_avalon_universal_slave_0_readdata
	wire         mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_waitrequest;     // traffic_controller_ch_8_9:uav_waitrequest -> mm_interconnect_1:traffic_controller_ch_8_9_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_debugaccess;     // mm_interconnect_1:traffic_controller_ch_8_9_avalon_universal_slave_0_debugaccess -> traffic_controller_ch_8_9:uav_debugaccess
	wire  [13:0] mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_address;         // mm_interconnect_1:traffic_controller_ch_8_9_avalon_universal_slave_0_address -> traffic_controller_ch_8_9:uav_address
	wire         mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_read;            // mm_interconnect_1:traffic_controller_ch_8_9_avalon_universal_slave_0_read -> traffic_controller_ch_8_9:uav_read
	wire   [3:0] mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_byteenable;      // mm_interconnect_1:traffic_controller_ch_8_9_avalon_universal_slave_0_byteenable -> traffic_controller_ch_8_9:uav_byteenable
	wire         mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_readdatavalid;   // traffic_controller_ch_8_9:uav_readdatavalid -> mm_interconnect_1:traffic_controller_ch_8_9_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_lock;            // mm_interconnect_1:traffic_controller_ch_8_9_avalon_universal_slave_0_lock -> traffic_controller_ch_8_9:uav_lock
	wire         mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_write;           // mm_interconnect_1:traffic_controller_ch_8_9_avalon_universal_slave_0_write -> traffic_controller_ch_8_9:uav_write
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_writedata;       // mm_interconnect_1:traffic_controller_ch_8_9_avalon_universal_slave_0_writedata -> traffic_controller_ch_8_9:uav_writedata
	wire   [2:0] mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_burstcount;      // mm_interconnect_1:traffic_controller_ch_8_9_avalon_universal_slave_0_burstcount -> traffic_controller_ch_8_9:uav_burstcount
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_readdata;      // traffic_controller_ch_10_11:uav_readdata -> mm_interconnect_1:traffic_controller_ch_10_11_avalon_universal_slave_0_readdata
	wire         mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_waitrequest;   // traffic_controller_ch_10_11:uav_waitrequest -> mm_interconnect_1:traffic_controller_ch_10_11_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_debugaccess;   // mm_interconnect_1:traffic_controller_ch_10_11_avalon_universal_slave_0_debugaccess -> traffic_controller_ch_10_11:uav_debugaccess
	wire  [13:0] mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_address;       // mm_interconnect_1:traffic_controller_ch_10_11_avalon_universal_slave_0_address -> traffic_controller_ch_10_11:uav_address
	wire         mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_read;          // mm_interconnect_1:traffic_controller_ch_10_11_avalon_universal_slave_0_read -> traffic_controller_ch_10_11:uav_read
	wire   [3:0] mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_byteenable;    // mm_interconnect_1:traffic_controller_ch_10_11_avalon_universal_slave_0_byteenable -> traffic_controller_ch_10_11:uav_byteenable
	wire         mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_readdatavalid; // traffic_controller_ch_10_11:uav_readdatavalid -> mm_interconnect_1:traffic_controller_ch_10_11_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_lock;          // mm_interconnect_1:traffic_controller_ch_10_11_avalon_universal_slave_0_lock -> traffic_controller_ch_10_11:uav_lock
	wire         mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_write;         // mm_interconnect_1:traffic_controller_ch_10_11_avalon_universal_slave_0_write -> traffic_controller_ch_10_11:uav_write
	wire  [31:0] mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_writedata;     // mm_interconnect_1:traffic_controller_ch_10_11_avalon_universal_slave_0_writedata -> traffic_controller_ch_10_11:uav_writedata
	wire   [2:0] mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_burstcount;    // mm_interconnect_1:traffic_controller_ch_10_11_avalon_universal_slave_0_burstcount -> traffic_controller_ch_10_11:uav_burstcount
	wire         rst_controller_reset_out_reset;                                                       // rst_controller:reset_out -> [master:reset, mm_clock_crossing_bridge:s0_reset, mm_interconnect_0:master_reset_reset_bridge_in_reset_reset, multi_channel:reset]
	wire         csr_clk_clk_reset_reset;                                                              // csr_clk:reset_n_out -> rst_controller:reset_in0
	wire         rst_controller_001_reset_out_reset;                                                   // rst_controller_001:reset_out -> [mm_clock_crossing_bridge:m0_reset, mm_interconnect_1:mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset, traffic_controller_ch_0_1:reset, traffic_controller_ch_10_11:reset, traffic_controller_ch_2_3:reset, traffic_controller_ch_4_5:reset, traffic_controller_ch_6_7:reset, traffic_controller_ch_8_9:reset]
	wire         mac_clk_clk_reset_reset;                                                              // mac_clk:reset_n_out -> rst_controller_001:reset_in0

	address_decoder_top_csr_clk csr_clk (
		.clk_out     (csr_clk_clk_clk),         //  output,  width = 1,          clk.clk
		.in_clk      (csr_clk_clk),             //   input,  width = 1,       clk_in.clk
		.reset_n     (csr_clk_reset_reset_n),   //   input,  width = 1, clk_in_reset.reset_n
		.reset_n_out (csr_clk_clk_reset_reset)  //  output,  width = 1,    clk_reset.reset_n
	);

	address_decoder_top_mac_clk mac_clk (
		.clk_out     (mac_clk_clk_clk),         //  output,  width = 1,          clk.clk
		.in_clk      (mac_clk_clk),             //   input,  width = 1,       clk_in.clk
		.reset_n     (mac_clk_reset_reset_n),   //   input,  width = 1, clk_in_reset.reset_n
		.reset_n_out (mac_clk_clk_reset_reset)  //  output,  width = 1,    clk_reset.reset_n
	);

	address_decoder_top_master master (
		.av_address        (slave_address),                                  //   input,  width = 26,      avalon_anti_master_0.address
		.av_waitrequest    (slave_waitrequest),                              //  output,   width = 1,                          .waitrequest
		.av_read           (slave_read),                                     //   input,   width = 1,                          .read
		.av_readdata       (slave_readdata),                                 //  output,  width = 32,                          .readdata
		.av_readdatavalid  (slave_readdatavalid),                            //  output,   width = 1,                          .readdatavalid
		.av_write          (slave_write),                                    //   input,   width = 1,                          .write
		.av_writedata      (slave_writedata),                                //   input,  width = 32,                          .writedata
		.uav_address       (master_avalon_universal_master_0_address),       //  output,  width = 32, avalon_universal_master_0.address
		.uav_burstcount    (master_avalon_universal_master_0_burstcount),    //  output,   width = 3,                          .burstcount
		.uav_read          (master_avalon_universal_master_0_read),          //  output,   width = 1,                          .read
		.uav_write         (master_avalon_universal_master_0_write),         //  output,   width = 1,                          .write
		.uav_waitrequest   (master_avalon_universal_master_0_waitrequest),   //   input,   width = 1,                          .waitrequest
		.uav_readdatavalid (master_avalon_universal_master_0_readdatavalid), //   input,   width = 1,                          .readdatavalid
		.uav_byteenable    (master_avalon_universal_master_0_byteenable),    //  output,   width = 4,                          .byteenable
		.uav_readdata      (master_avalon_universal_master_0_readdata),      //   input,  width = 32,                          .readdata
		.uav_writedata     (master_avalon_universal_master_0_writedata),     //  output,  width = 32,                          .writedata
		.uav_lock          (master_avalon_universal_master_0_lock),          //  output,   width = 1,                          .lock
		.uav_debugaccess   (master_avalon_universal_master_0_debugaccess),   //  output,   width = 1,                          .debugaccess
		.clk               (csr_clk_clk_clk),                                //   input,   width = 1,                       clk.clk
		.reset             (rst_controller_reset_out_reset)                  //   input,   width = 1,                     reset.reset
	);

	address_decoder_top_mm_clock_crossing_bridge mm_clock_crossing_bridge (
		.m0_waitrequest   (mm_clock_crossing_bridge_m0_waitrequest),                     //   input,   width = 1,       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_m0_readdata),                        //   input,  width = 32,         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_m0_readdatavalid),                   //   input,   width = 1,         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_m0_burstcount),                      //  output,   width = 1,         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_m0_writedata),                       //  output,  width = 32,         .writedata
		.m0_address       (mm_clock_crossing_bridge_m0_address),                         //  output,  width = 17,         .address
		.m0_write         (mm_clock_crossing_bridge_m0_write),                           //  output,   width = 1,         .write
		.m0_read          (mm_clock_crossing_bridge_m0_read),                            //  output,   width = 1,         .read
		.m0_byteenable    (mm_clock_crossing_bridge_m0_byteenable),                      //  output,   width = 4,         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_m0_debugaccess),                     //  output,   width = 1,         .debugaccess
		.m0_clk           (mac_clk_clk_clk),                                             //   input,   width = 1,   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                          //   input,   width = 1, m0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),   //  output,   width = 1,       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),      //  output,  width = 32,         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid), //  output,   width = 1,         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),    //   input,   width = 1,         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),     //   input,  width = 32,         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),       //   input,  width = 17,         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),         //   input,   width = 1,         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),          //   input,   width = 1,         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),    //   input,   width = 4,         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),   //   input,   width = 1,         .debugaccess
		.s0_clk           (csr_clk_clk_clk),                                             //   input,   width = 1,   s0_clk.clk
		.s0_reset         (rst_controller_reset_out_reset)                               //   input,   width = 1, s0_reset.reset
	);

	address_decoder_top_multi_channel multi_channel (
		.av_address        (multi_channel_address),                                                  //  output,  width = 20,      avalon_anti_slave_0.address
		.av_write          (multi_channel_write),                                                    //  output,   width = 1,                         .write
		.av_read           (multi_channel_read),                                                     //  output,   width = 1,                         .read
		.av_readdata       (multi_channel_readdata),                                                 //   input,  width = 32,                         .readdata
		.av_writedata      (multi_channel_writedata),                                                //  output,  width = 32,                         .writedata
		.av_waitrequest    (multi_channel_waitrequest),                                              //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_multi_channel_avalon_universal_slave_0_address),       //   input,  width = 20, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_multi_channel_avalon_universal_slave_0_burstcount),    //   input,   width = 3,                         .burstcount
		.uav_read          (mm_interconnect_0_multi_channel_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_multi_channel_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_multi_channel_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_multi_channel_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_multi_channel_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_multi_channel_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_multi_channel_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_multi_channel_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_multi_channel_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (csr_clk_clk_clk),                                                        //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decoder_top_traffic_controller_ch_0_1 traffic_controller_ch_0_1 (
		.av_address        (traffic_controller_ch_0_1_address),                                                  //  output,  width = 14,      avalon_anti_slave_0.address
		.av_write          (traffic_controller_ch_0_1_write),                                                    //  output,   width = 1,                         .write
		.av_read           (traffic_controller_ch_0_1_read),                                                     //  output,   width = 1,                         .read
		.av_readdata       (traffic_controller_ch_0_1_readdata),                                                 //   input,  width = 32,                         .readdata
		.av_writedata      (traffic_controller_ch_0_1_writedata),                                                //  output,  width = 32,                         .writedata
		.av_waitrequest    (traffic_controller_ch_0_1_waitrequest),                                              //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_burstcount),    //   input,   width = 3,                         .burstcount
		.uav_read          (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (mac_clk_clk_clk),                                                                    //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_001_reset_out_reset)                                                  //   input,   width = 1,                    reset.reset
	);

	address_decoder_top_traffic_controller_ch_10_11 traffic_controller_ch_10_11 (
		.av_address        (traffic_controller_ch_10_11_address),                                                  //  output,  width = 14,      avalon_anti_slave_0.address
		.av_write          (traffic_controller_ch_10_11_write),                                                    //  output,   width = 1,                         .write
		.av_read           (traffic_controller_ch_10_11_read),                                                     //  output,   width = 1,                         .read
		.av_readdata       (traffic_controller_ch_10_11_readdata),                                                 //   input,  width = 32,                         .readdata
		.av_writedata      (traffic_controller_ch_10_11_writedata),                                                //  output,  width = 32,                         .writedata
		.av_waitrequest    (traffic_controller_ch_10_11_waitrequest),                                              //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_burstcount),    //   input,   width = 3,                         .burstcount
		.uav_read          (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (mac_clk_clk_clk),                                                                      //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_001_reset_out_reset)                                                    //   input,   width = 1,                    reset.reset
	);

	address_decoder_top_traffic_controller_ch_2_3 traffic_controller_ch_2_3 (
		.av_address        (traffic_controller_ch_2_3_address),                                                  //  output,  width = 14,      avalon_anti_slave_0.address
		.av_write          (traffic_controller_ch_2_3_write),                                                    //  output,   width = 1,                         .write
		.av_read           (traffic_controller_ch_2_3_read),                                                     //  output,   width = 1,                         .read
		.av_readdata       (traffic_controller_ch_2_3_readdata),                                                 //   input,  width = 32,                         .readdata
		.av_writedata      (traffic_controller_ch_2_3_writedata),                                                //  output,  width = 32,                         .writedata
		.av_waitrequest    (traffic_controller_ch_2_3_waitrequest),                                              //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_burstcount),    //   input,   width = 3,                         .burstcount
		.uav_read          (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (mac_clk_clk_clk),                                                                    //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_001_reset_out_reset)                                                  //   input,   width = 1,                    reset.reset
	);

	address_decoder_top_traffic_controller_ch_4_5 traffic_controller_ch_4_5 (
		.av_address        (traffic_controller_ch_4_5_address),                                                  //  output,  width = 14,      avalon_anti_slave_0.address
		.av_write          (traffic_controller_ch_4_5_write),                                                    //  output,   width = 1,                         .write
		.av_read           (traffic_controller_ch_4_5_read),                                                     //  output,   width = 1,                         .read
		.av_readdata       (traffic_controller_ch_4_5_readdata),                                                 //   input,  width = 32,                         .readdata
		.av_writedata      (traffic_controller_ch_4_5_writedata),                                                //  output,  width = 32,                         .writedata
		.av_waitrequest    (traffic_controller_ch_4_5_waitrequest),                                              //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_burstcount),    //   input,   width = 3,                         .burstcount
		.uav_read          (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (mac_clk_clk_clk),                                                                    //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_001_reset_out_reset)                                                  //   input,   width = 1,                    reset.reset
	);

	address_decoder_top_traffic_controller_ch_6_7 traffic_controller_ch_6_7 (
		.av_address        (traffic_controller_ch_6_7_address),                                                  //  output,  width = 14,      avalon_anti_slave_0.address
		.av_write          (traffic_controller_ch_6_7_write),                                                    //  output,   width = 1,                         .write
		.av_read           (traffic_controller_ch_6_7_read),                                                     //  output,   width = 1,                         .read
		.av_readdata       (traffic_controller_ch_6_7_readdata),                                                 //   input,  width = 32,                         .readdata
		.av_writedata      (traffic_controller_ch_6_7_writedata),                                                //  output,  width = 32,                         .writedata
		.av_waitrequest    (traffic_controller_ch_6_7_waitrequest),                                              //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_burstcount),    //   input,   width = 3,                         .burstcount
		.uav_read          (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (mac_clk_clk_clk),                                                                    //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_001_reset_out_reset)                                                  //   input,   width = 1,                    reset.reset
	);

	address_decoder_top_traffic_controller_ch_8_9 traffic_controller_ch_8_9 (
		.av_address        (traffic_controller_ch_8_9_address),                                                  //  output,  width = 14,      avalon_anti_slave_0.address
		.av_write          (traffic_controller_ch_8_9_write),                                                    //  output,   width = 1,                         .write
		.av_read           (traffic_controller_ch_8_9_read),                                                     //  output,   width = 1,                         .read
		.av_readdata       (traffic_controller_ch_8_9_readdata),                                                 //   input,  width = 32,                         .readdata
		.av_writedata      (traffic_controller_ch_8_9_writedata),                                                //  output,  width = 32,                         .writedata
		.av_waitrequest    (traffic_controller_ch_8_9_waitrequest),                                              //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_burstcount),    //   input,   width = 3,                         .burstcount
		.uav_read          (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (mac_clk_clk_clk),                                                                    //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_001_reset_out_reset)                                                  //   input,   width = 1,                    reset.reset
	);

	address_decoder_top_altera_mm_interconnect_1920_tgojdoy mm_interconnect_0 (
		.master_avalon_universal_master_0_address             (master_avalon_universal_master_0_address),                               //   input,  width = 32,       master_avalon_universal_master_0.address
		.master_avalon_universal_master_0_waitrequest         (master_avalon_universal_master_0_waitrequest),                           //  output,   width = 1,                                       .waitrequest
		.master_avalon_universal_master_0_burstcount          (master_avalon_universal_master_0_burstcount),                            //   input,   width = 3,                                       .burstcount
		.master_avalon_universal_master_0_byteenable          (master_avalon_universal_master_0_byteenable),                            //   input,   width = 4,                                       .byteenable
		.master_avalon_universal_master_0_read                (master_avalon_universal_master_0_read),                                  //   input,   width = 1,                                       .read
		.master_avalon_universal_master_0_readdata            (master_avalon_universal_master_0_readdata),                              //  output,  width = 32,                                       .readdata
		.master_avalon_universal_master_0_readdatavalid       (master_avalon_universal_master_0_readdatavalid),                         //  output,   width = 1,                                       .readdatavalid
		.master_avalon_universal_master_0_write               (master_avalon_universal_master_0_write),                                 //   input,   width = 1,                                       .write
		.master_avalon_universal_master_0_writedata           (master_avalon_universal_master_0_writedata),                             //   input,  width = 32,                                       .writedata
		.master_avalon_universal_master_0_lock                (master_avalon_universal_master_0_lock),                                  //   input,   width = 1,                                       .lock
		.master_avalon_universal_master_0_debugaccess         (master_avalon_universal_master_0_debugaccess),                           //   input,   width = 1,                                       .debugaccess
		.multi_channel_avalon_universal_slave_0_address       (mm_interconnect_0_multi_channel_avalon_universal_slave_0_address),       //  output,  width = 20, multi_channel_avalon_universal_slave_0.address
		.multi_channel_avalon_universal_slave_0_write         (mm_interconnect_0_multi_channel_avalon_universal_slave_0_write),         //  output,   width = 1,                                       .write
		.multi_channel_avalon_universal_slave_0_read          (mm_interconnect_0_multi_channel_avalon_universal_slave_0_read),          //  output,   width = 1,                                       .read
		.multi_channel_avalon_universal_slave_0_readdata      (mm_interconnect_0_multi_channel_avalon_universal_slave_0_readdata),      //   input,  width = 32,                                       .readdata
		.multi_channel_avalon_universal_slave_0_writedata     (mm_interconnect_0_multi_channel_avalon_universal_slave_0_writedata),     //  output,  width = 32,                                       .writedata
		.multi_channel_avalon_universal_slave_0_burstcount    (mm_interconnect_0_multi_channel_avalon_universal_slave_0_burstcount),    //  output,   width = 3,                                       .burstcount
		.multi_channel_avalon_universal_slave_0_byteenable    (mm_interconnect_0_multi_channel_avalon_universal_slave_0_byteenable),    //  output,   width = 4,                                       .byteenable
		.multi_channel_avalon_universal_slave_0_readdatavalid (mm_interconnect_0_multi_channel_avalon_universal_slave_0_readdatavalid), //   input,   width = 1,                                       .readdatavalid
		.multi_channel_avalon_universal_slave_0_waitrequest   (mm_interconnect_0_multi_channel_avalon_universal_slave_0_waitrequest),   //   input,   width = 1,                                       .waitrequest
		.multi_channel_avalon_universal_slave_0_lock          (mm_interconnect_0_multi_channel_avalon_universal_slave_0_lock),          //  output,   width = 1,                                       .lock
		.multi_channel_avalon_universal_slave_0_debugaccess   (mm_interconnect_0_multi_channel_avalon_universal_slave_0_debugaccess),   //  output,   width = 1,                                       .debugaccess
		.mm_clock_crossing_bridge_s0_address                  (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),                  //  output,  width = 17,            mm_clock_crossing_bridge_s0.address
		.mm_clock_crossing_bridge_s0_write                    (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),                    //  output,   width = 1,                                       .write
		.mm_clock_crossing_bridge_s0_read                     (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),                     //  output,   width = 1,                                       .read
		.mm_clock_crossing_bridge_s0_readdata                 (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),                 //   input,  width = 32,                                       .readdata
		.mm_clock_crossing_bridge_s0_writedata                (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),                //  output,  width = 32,                                       .writedata
		.mm_clock_crossing_bridge_s0_burstcount               (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),               //  output,   width = 1,                                       .burstcount
		.mm_clock_crossing_bridge_s0_byteenable               (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),               //  output,   width = 4,                                       .byteenable
		.mm_clock_crossing_bridge_s0_readdatavalid            (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid),            //   input,   width = 1,                                       .readdatavalid
		.mm_clock_crossing_bridge_s0_waitrequest              (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),              //   input,   width = 1,                                       .waitrequest
		.mm_clock_crossing_bridge_s0_debugaccess              (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),              //  output,   width = 1,                                       .debugaccess
		.master_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                                         //   input,   width = 1,     master_reset_reset_bridge_in_reset.reset
		.csr_clk_clk_clk                                      (csr_clk_clk_clk)                                                         //   input,   width = 1,                            csr_clk_clk.clk
	);

	address_decoder_top_altera_mm_interconnect_1920_4grhzia mm_interconnect_1 (
		.mm_clock_crossing_bridge_m0_address                                (mm_clock_crossing_bridge_m0_address),                                                  //   input,  width = 17,                             mm_clock_crossing_bridge_m0.address
		.mm_clock_crossing_bridge_m0_waitrequest                            (mm_clock_crossing_bridge_m0_waitrequest),                                              //  output,   width = 1,                                                        .waitrequest
		.mm_clock_crossing_bridge_m0_burstcount                             (mm_clock_crossing_bridge_m0_burstcount),                                               //   input,   width = 1,                                                        .burstcount
		.mm_clock_crossing_bridge_m0_byteenable                             (mm_clock_crossing_bridge_m0_byteenable),                                               //   input,   width = 4,                                                        .byteenable
		.mm_clock_crossing_bridge_m0_read                                   (mm_clock_crossing_bridge_m0_read),                                                     //   input,   width = 1,                                                        .read
		.mm_clock_crossing_bridge_m0_readdata                               (mm_clock_crossing_bridge_m0_readdata),                                                 //  output,  width = 32,                                                        .readdata
		.mm_clock_crossing_bridge_m0_readdatavalid                          (mm_clock_crossing_bridge_m0_readdatavalid),                                            //  output,   width = 1,                                                        .readdatavalid
		.mm_clock_crossing_bridge_m0_write                                  (mm_clock_crossing_bridge_m0_write),                                                    //   input,   width = 1,                                                        .write
		.mm_clock_crossing_bridge_m0_writedata                              (mm_clock_crossing_bridge_m0_writedata),                                                //   input,  width = 32,                                                        .writedata
		.mm_clock_crossing_bridge_m0_debugaccess                            (mm_clock_crossing_bridge_m0_debugaccess),                                              //   input,   width = 1,                                                        .debugaccess
		.traffic_controller_ch_0_1_avalon_universal_slave_0_address         (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_address),         //  output,  width = 14,      traffic_controller_ch_0_1_avalon_universal_slave_0.address
		.traffic_controller_ch_0_1_avalon_universal_slave_0_write           (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_write),           //  output,   width = 1,                                                        .write
		.traffic_controller_ch_0_1_avalon_universal_slave_0_read            (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_read),            //  output,   width = 1,                                                        .read
		.traffic_controller_ch_0_1_avalon_universal_slave_0_readdata        (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                        .readdata
		.traffic_controller_ch_0_1_avalon_universal_slave_0_writedata       (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                        .writedata
		.traffic_controller_ch_0_1_avalon_universal_slave_0_burstcount      (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_burstcount),      //  output,   width = 3,                                                        .burstcount
		.traffic_controller_ch_0_1_avalon_universal_slave_0_byteenable      (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                        .byteenable
		.traffic_controller_ch_0_1_avalon_universal_slave_0_readdatavalid   (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                        .readdatavalid
		.traffic_controller_ch_0_1_avalon_universal_slave_0_waitrequest     (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                        .waitrequest
		.traffic_controller_ch_0_1_avalon_universal_slave_0_lock            (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                        .lock
		.traffic_controller_ch_0_1_avalon_universal_slave_0_debugaccess     (mm_interconnect_1_traffic_controller_ch_0_1_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                        .debugaccess
		.traffic_controller_ch_2_3_avalon_universal_slave_0_address         (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_address),         //  output,  width = 14,      traffic_controller_ch_2_3_avalon_universal_slave_0.address
		.traffic_controller_ch_2_3_avalon_universal_slave_0_write           (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_write),           //  output,   width = 1,                                                        .write
		.traffic_controller_ch_2_3_avalon_universal_slave_0_read            (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_read),            //  output,   width = 1,                                                        .read
		.traffic_controller_ch_2_3_avalon_universal_slave_0_readdata        (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                        .readdata
		.traffic_controller_ch_2_3_avalon_universal_slave_0_writedata       (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                        .writedata
		.traffic_controller_ch_2_3_avalon_universal_slave_0_burstcount      (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_burstcount),      //  output,   width = 3,                                                        .burstcount
		.traffic_controller_ch_2_3_avalon_universal_slave_0_byteenable      (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                        .byteenable
		.traffic_controller_ch_2_3_avalon_universal_slave_0_readdatavalid   (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                        .readdatavalid
		.traffic_controller_ch_2_3_avalon_universal_slave_0_waitrequest     (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                        .waitrequest
		.traffic_controller_ch_2_3_avalon_universal_slave_0_lock            (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                        .lock
		.traffic_controller_ch_2_3_avalon_universal_slave_0_debugaccess     (mm_interconnect_1_traffic_controller_ch_2_3_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                        .debugaccess
		.traffic_controller_ch_4_5_avalon_universal_slave_0_address         (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_address),         //  output,  width = 14,      traffic_controller_ch_4_5_avalon_universal_slave_0.address
		.traffic_controller_ch_4_5_avalon_universal_slave_0_write           (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_write),           //  output,   width = 1,                                                        .write
		.traffic_controller_ch_4_5_avalon_universal_slave_0_read            (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_read),            //  output,   width = 1,                                                        .read
		.traffic_controller_ch_4_5_avalon_universal_slave_0_readdata        (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                        .readdata
		.traffic_controller_ch_4_5_avalon_universal_slave_0_writedata       (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                        .writedata
		.traffic_controller_ch_4_5_avalon_universal_slave_0_burstcount      (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_burstcount),      //  output,   width = 3,                                                        .burstcount
		.traffic_controller_ch_4_5_avalon_universal_slave_0_byteenable      (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                        .byteenable
		.traffic_controller_ch_4_5_avalon_universal_slave_0_readdatavalid   (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                        .readdatavalid
		.traffic_controller_ch_4_5_avalon_universal_slave_0_waitrequest     (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                        .waitrequest
		.traffic_controller_ch_4_5_avalon_universal_slave_0_lock            (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                        .lock
		.traffic_controller_ch_4_5_avalon_universal_slave_0_debugaccess     (mm_interconnect_1_traffic_controller_ch_4_5_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                        .debugaccess
		.traffic_controller_ch_6_7_avalon_universal_slave_0_address         (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_address),         //  output,  width = 14,      traffic_controller_ch_6_7_avalon_universal_slave_0.address
		.traffic_controller_ch_6_7_avalon_universal_slave_0_write           (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_write),           //  output,   width = 1,                                                        .write
		.traffic_controller_ch_6_7_avalon_universal_slave_0_read            (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_read),            //  output,   width = 1,                                                        .read
		.traffic_controller_ch_6_7_avalon_universal_slave_0_readdata        (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                        .readdata
		.traffic_controller_ch_6_7_avalon_universal_slave_0_writedata       (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                        .writedata
		.traffic_controller_ch_6_7_avalon_universal_slave_0_burstcount      (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_burstcount),      //  output,   width = 3,                                                        .burstcount
		.traffic_controller_ch_6_7_avalon_universal_slave_0_byteenable      (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                        .byteenable
		.traffic_controller_ch_6_7_avalon_universal_slave_0_readdatavalid   (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                        .readdatavalid
		.traffic_controller_ch_6_7_avalon_universal_slave_0_waitrequest     (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                        .waitrequest
		.traffic_controller_ch_6_7_avalon_universal_slave_0_lock            (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                        .lock
		.traffic_controller_ch_6_7_avalon_universal_slave_0_debugaccess     (mm_interconnect_1_traffic_controller_ch_6_7_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                        .debugaccess
		.traffic_controller_ch_8_9_avalon_universal_slave_0_address         (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_address),         //  output,  width = 14,      traffic_controller_ch_8_9_avalon_universal_slave_0.address
		.traffic_controller_ch_8_9_avalon_universal_slave_0_write           (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_write),           //  output,   width = 1,                                                        .write
		.traffic_controller_ch_8_9_avalon_universal_slave_0_read            (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_read),            //  output,   width = 1,                                                        .read
		.traffic_controller_ch_8_9_avalon_universal_slave_0_readdata        (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                        .readdata
		.traffic_controller_ch_8_9_avalon_universal_slave_0_writedata       (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                        .writedata
		.traffic_controller_ch_8_9_avalon_universal_slave_0_burstcount      (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_burstcount),      //  output,   width = 3,                                                        .burstcount
		.traffic_controller_ch_8_9_avalon_universal_slave_0_byteenable      (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                        .byteenable
		.traffic_controller_ch_8_9_avalon_universal_slave_0_readdatavalid   (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                        .readdatavalid
		.traffic_controller_ch_8_9_avalon_universal_slave_0_waitrequest     (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                        .waitrequest
		.traffic_controller_ch_8_9_avalon_universal_slave_0_lock            (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                        .lock
		.traffic_controller_ch_8_9_avalon_universal_slave_0_debugaccess     (mm_interconnect_1_traffic_controller_ch_8_9_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                        .debugaccess
		.traffic_controller_ch_10_11_avalon_universal_slave_0_address       (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_address),       //  output,  width = 14,    traffic_controller_ch_10_11_avalon_universal_slave_0.address
		.traffic_controller_ch_10_11_avalon_universal_slave_0_write         (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_write),         //  output,   width = 1,                                                        .write
		.traffic_controller_ch_10_11_avalon_universal_slave_0_read          (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_read),          //  output,   width = 1,                                                        .read
		.traffic_controller_ch_10_11_avalon_universal_slave_0_readdata      (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_readdata),      //   input,  width = 32,                                                        .readdata
		.traffic_controller_ch_10_11_avalon_universal_slave_0_writedata     (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_writedata),     //  output,  width = 32,                                                        .writedata
		.traffic_controller_ch_10_11_avalon_universal_slave_0_burstcount    (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_burstcount),    //  output,   width = 3,                                                        .burstcount
		.traffic_controller_ch_10_11_avalon_universal_slave_0_byteenable    (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_byteenable),    //  output,   width = 4,                                                        .byteenable
		.traffic_controller_ch_10_11_avalon_universal_slave_0_readdatavalid (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_readdatavalid), //   input,   width = 1,                                                        .readdatavalid
		.traffic_controller_ch_10_11_avalon_universal_slave_0_waitrequest   (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_waitrequest),   //   input,   width = 1,                                                        .waitrequest
		.traffic_controller_ch_10_11_avalon_universal_slave_0_lock          (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_lock),          //  output,   width = 1,                                                        .lock
		.traffic_controller_ch_10_11_avalon_universal_slave_0_debugaccess   (mm_interconnect_1_traffic_controller_ch_10_11_avalon_universal_slave_0_debugaccess),   //  output,   width = 1,                                                        .debugaccess
		.mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                                                   //   input,   width = 1, mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset.reset
		.mac_clk_clk_clk                                                    (mac_clk_clk_clk)                                                                       //   input,   width = 1,                                             mac_clk_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~csr_clk_clk_reset_reset),       //   input,  width = 1, reset_in0.reset
		.clk            (csr_clk_clk_clk),                //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                               // (terminated),                       
		.reset_req_in0  (1'b0),                           // (terminated),                       
		.reset_in1      (1'b0),                           // (terminated),                       
		.reset_req_in1  (1'b0),                           // (terminated),                       
		.reset_in2      (1'b0),                           // (terminated),                       
		.reset_req_in2  (1'b0),                           // (terminated),                       
		.reset_in3      (1'b0),                           // (terminated),                       
		.reset_req_in3  (1'b0),                           // (terminated),                       
		.reset_in4      (1'b0),                           // (terminated),                       
		.reset_req_in4  (1'b0),                           // (terminated),                       
		.reset_in5      (1'b0),                           // (terminated),                       
		.reset_req_in5  (1'b0),                           // (terminated),                       
		.reset_in6      (1'b0),                           // (terminated),                       
		.reset_req_in6  (1'b0),                           // (terminated),                       
		.reset_in7      (1'b0),                           // (terminated),                       
		.reset_req_in7  (1'b0),                           // (terminated),                       
		.reset_in8      (1'b0),                           // (terminated),                       
		.reset_req_in8  (1'b0),                           // (terminated),                       
		.reset_in9      (1'b0),                           // (terminated),                       
		.reset_req_in9  (1'b0),                           // (terminated),                       
		.reset_in10     (1'b0),                           // (terminated),                       
		.reset_req_in10 (1'b0),                           // (terminated),                       
		.reset_in11     (1'b0),                           // (terminated),                       
		.reset_req_in11 (1'b0),                           // (terminated),                       
		.reset_in12     (1'b0),                           // (terminated),                       
		.reset_req_in12 (1'b0),                           // (terminated),                       
		.reset_in13     (1'b0),                           // (terminated),                       
		.reset_req_in13 (1'b0),                           // (terminated),                       
		.reset_in14     (1'b0),                           // (terminated),                       
		.reset_req_in14 (1'b0),                           // (terminated),                       
		.reset_in15     (1'b0),                           // (terminated),                       
		.reset_req_in15 (1'b0)                            // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~mac_clk_clk_reset_reset),           //   input,  width = 1, reset_in0.reset
		.clk            (mac_clk_clk_clk),                    //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
