// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
g3nCyV1P1iaIGYvOr2BuE8X6K6HQ1rb6YCaxjnRV39hDQtGcltRWzFIfU9za
TC1SoEsFZui1vjkAs9JtmJ7eKxz1l5TouzdKHmGj8SbSfq9YbhVezkxGwPo5
iSvna0nskbu2X4c740jjCdWBFvg+zZq1IJMhRyG3HKsgpWikfLkguUnRK3gA
CDXFaU6CY+Tpm/6dQJFKVE32t7o9xhlEg6RiTJvzs/ehtLDRqf289DdsCHxK
YfWmxW08yISG1bgvUEESmsXkqmG+ETVTDg69o2rdcVeNCAhzaAsLtQjfxYhR
U38ynqlD1OgQ9cizepNEvRCf/ZhwDqpw/SlG7i72Vw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CwxdaFNhGXdNPQ6j7TJ/clwDWNYp4cIMZkW7EJ4vPmVV6GPHFTMefSRNyIci
VJ4WQj3+g/XatmdAiwFV3Y2hF4t/WzbNtSjKy9Q+ivpSARXuC4sxkJ3O9BMh
dH0X3SruDn4LbzjJxuvOEAl13Uhxdt9RLt3lNf8IXGJSFgQ0A5XL0nHtVzZK
XSRz85gKduGghC6JqYSSJNijmitMc2JgbeMU3hzJ/riz/V01vlW1iRmCdCa9
mbas0qlJEzRPFR8eVNSmhoDFwttsaUIFoevCEBsuZk12ytXBxxNfyEp1Usfx
bHYi9jRCdSxg+fHSs251oqTjJ6SYFNDTWPBJgrDdlg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Y+kuvR5QQ0GwrYMymTqLmUZ2lLJi3/766iCLlYC6y4uzc0Y9wkaLq4RjHcAi
h8dg1RYxZ4wGwwXd01Cf+Jzp/Vj1YCmnLiaOe+y4RXlB0JipkGOQtMQga6tM
37iQpR4YxsSc2cTjYcCf/Ea4lr+r0kRsu2VbzKLd5DYv7WOriLtRmDvQ7oRm
witW1oxzDTxH8Qk9il1dg8gefq2rQD571CO1FjMlvkv5HCaar/63ZZIegsmf
IlrorJErPFLO74gimjyCSg38xizOCOFvLMybG1j8Zu/2JPbm65sHeYkh+z7n
EtsnHYQbEhy3DuyreeKNGzY+n4G357awshFci3ZVSQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
g8Rkq50HzFH28Vr609OQY/UTvmhve69WiKR9+KOVtNXlNeT4H5UYlKW5PKDx
Afh02aKts2k2ye8h/0+Xryk2xP/2FfmtdrC33qcqSbcMoDJgob0jTk9Gh8wV
XkQv6e/PQAKSkUHi33wRkVYremOLFPcaaLibZZpzKTFI9a0V9pU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NCdfd8aHY2grXzjKRgkxVMenVhADrlhDGqUIfZW3Nse+vjNTsJfvGGSdUvcm
ZjHUqe0JPWggeO+4xG+YmyGTXarUS4+2/Rpy8gyPpBd9zbBw/OBf0+f+3gXv
6dltj/3YdBbueHFnjo5tOkYnN6wv0na74U09G8zIx0CIJzAxTtb8em9q6wvI
V6J6f6wNZUd1juAweLkkNGtnvfXQuOEYflclt07gyOHAGuosInVS0sgiCotq
+Rl9BGwx1zRIwG1MQ7GS1yBfYCGv7Pgwr6c7jegm52uswJSaAoBBQJLOUvfD
0PxnH4YrUGw1niCyX9utXOpYdNcaq1ULaXdRs4MJHOLhdX8We7EVfJRKHWDw
H/SWKYYOH6Hc+R+va86JY+yGPBRGB989rClCxxI+mHPRh+jhkawC3/jYMMY+
l7nMFcPvfg1ykyyyF7WZQRIAfTy5FpJQpU1912PIVu0xQnwWfhkr6foFVtgK
yiPPzceIcr8iFNn1xDh+5eusLDcS2eB7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A7YcsX4EyfzQ+mC1XBMzKVAqxqJtwXkYNPopvmzOcw1NODhB+88Px43S6nE/
T014yW7YEqeMlBveNOZoGEY3Si0DkVtU6KGxSAVgHF5k/y8FOzjFsvUkkjr+
xWkTxtJW7YfpqYBx6+yG4xipwBizZ3Fe1W8Si4XL1lU/bZazadQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PFWjaMHzpp56PDRd+RSWlQ0yTfWy/Dmr1MFFN82O9ssZ3qfOKBgE70vio666
sHp+Ym8QW2f1FTst32QghdNWkh9PVsL5qy5OnOrXVPret2gE9ij+slDR4pPm
C+j5ay+tZDQWuEohxAlq0PvcysVU8KSpcJkSZ9hFgIhYYv6/KKg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 91312)
`pragma protect data_block
1quG+JN9lMtalNZw7ysFdWzS9ACQKWlADkIa/lwvLrGB+dxAOL66XtpcvEWQ
1g1lqIlu3npPDepTPTGGKW5fjftKTCVQn0rzCrk5nj0/OvGIOjnbExbHJBXO
QLP750tIJZA5C1EWd9gsg8T60/b/Xk+5HvALbk6kbdl/nn2JM4mNZolrdtVF
Me6OqoOGEabkeOF5Z4yewtP3J0UwZLViPsDwzIlKLUWRgdu4n22j8KOl7+8Y
V6sIei2jUkRT2lEYIEvafA3iWwV+d5uBF8ti0vzith9L/POiFMmGD+Mb6+vP
rSyN9KiEapPc8jLeO0HsqCiQigOcoS9Mx2g1GF01OLObhSfvHDmbJqrDwOqj
cfhYbG08VVdC5cHAw3FI3SczHKmt8X+osAnbgFV3TPP5B2hAgcWt/yHI0+rZ
ouGHPUoHWV3+ssC9UNw1DbvOfept0T5F5wzZh72/0wPdYA3+9vJ0dKzICIU2
OxFY98dnRzsnW+ODalS2ztOQTQfXRrvF6oAepl4J1aCMdaOPvkravKaIEtJ1
h5drRYjylpZQ2sTEgULCLfw91hopPPaMZ+QpKB/9pAG7Y1CNKOihdaLA84ys
+hOSVQdhdfi84wZiXltzufCBEQ7BV2Y3uX+agkydTaxon+qTE1tGg37P9MIE
QBOF/Q24QyyDvS/w4LQo+vUEkIXR2ltsqG1NBs0l0+07KJybvxhQQ40F+0uj
YdfoqSPAPzqgh61wSzcSDwCmyUJ8vcX2NNT4Fg9LV4gOxwJ9ZXHaXrB1XtSK
FaSl0Qgrqz0Iq930qzKkmhHIMhloA7MT8XaaXxTtUjU9pUp6OkeVrtboqv/P
JF9IRN+CwP90/QBq46frGhjeX7bq8ZV8ZBcJs8jzw0jscAmuSnVPex01+jT0
HeBcYcfbx0I4rlk7piIoltyMSBJ4QO+TzRxtTVrxf729wPEU1DOHmfIirdTN
TbeLVZ0OpAvvyAEQ3OzqaKMyL7ZmzLbRb73GigbJQmEgnEkKM7LerckPxFkh
+Dzg60030ob9gCgM7MB0jiDVyQsSZCBh3rCKm1f2OqU39CdZSg0QZV+/e53P
CTjnuq2eUnlsdXIOV/+3KtpfZKWeDv5qprJiGOP+mA9OeyyfY057Hvn1tISM
IxgdlIZQkjkdXg3Th7SCIRzqdx2Dzj+y17yjlYX66WRVJ0TXJPjPAxoMN6LI
qIMW/PcjQ+QP+cBFwv+NkJC338Fp7sU6JvbuO/MljgVFr+3k1WsI89iZiLdN
Gsu98j1un0OvXc3n2WZMC7hGuEZT5gXmpvObm1xS6U1vn3xiFcUMBbXMPlPq
TqAbu0kSg+IGSMLU3Q2gDhGsLw8c4TgnkGNLZxd1eHqUyBXeqtKOx4//dzhN
ZiUVYdcILrn5pMA7HemQbcPsykhSJTCtT7xeotJH9M9iBao2pqnMFcfUc7fN
nKhLD75CR9xYxMsqxLbYoIfmNrBYkZKpBfpJp2o7facDCAuL8crGqH+h99xI
N0Ugs4Rn8396Doyy7K02RaGLN4Pl7Qi3XAsAgUR4WWqhcCi1aBZUraKhh5iW
rSZamQFeqmyd0p4pxYAVQypmExQspRreZ11TIqg5J+Rsr9Lnboz8rRJqSyQk
dceQPEbMKLaqdT4vQTsUSalJGh0DGoXFEGPsO2ye7X9/CkEML4YSIS9ogKY1
wSTSjMiys+gNGkCfHKZywk5qdaYltcVx9kdsE0wCEm8kZQqJgEG+p0IThwrV
WBrO2Ya0+dTRTkaJZAzI4Jmo5GWPA1DeDH4E0tPfGE2uzs2DUCJosICHaCVZ
y/3QolGo1OBeCeszWgl0otj1b2iLxppLieIsB94etsBtC6Qp2mwh5aBk3IRh
rTonPdvj35ItVgQeWG+Uyeyhis63iMRKx+ukRB6wj3FzFh3IbQQ3TmYgGsc9
0vfX4ccxT72hcdyTMb9Lp++OCGrrsT+LQpiLv+kvdyonmiXt2+5GlpIy46t1
x6qj+SKnV+g2K49TmGw21VI66uaBsolr5cpIDSbXu9EMjhu9PXPecH69Hu+0
uoAyEFwUJo82G41KmmDmJnCMEHhEOvFJROd84eIuABfBLjhsSvC8VhWY6L4V
WkIrWAiwn1bMViYfx6E51PYbniYxarUfFPwC7cI4Y9OdoFnL2L3R15zVQonT
gmLLFGdEd611dAkguHyhF0xq9jL0euRPnnT5TpZjgIKUdsHyWm/qrS5kxSHf
hvaqc1w08+UYwnnCS+Rznr73XQwO1VQjT52QQu+bCIskf4hwZGabnuu56fB2
iOxhXWbj//iHlRGFbIeHXu9X+kfb7DZ2u5bSUVBxzS6b56YRRQkqicn22VBl
gT0jmfjEXRh836et1xCsPXU6wuLPnseOg+MvNHSWY/v24RKjqMZp79pjyyjj
/N79BsJPLa6FfmdG/U1B03OfUkrOX+WfiSvquQwq8FzaQs+O8DKtGyFISkSM
sT61Jpq3A/ZAfEqEAR+fX+in2HFRYR5sshh92FLRKke5WzMc9pGb4BrUCeeP
sAMSDPmHwEXxIOa1vloTMxZ7NEwCPmDNWLrPoHyJ+Ku4dAbGKJLn6BBUNFfd
SYpOTywe0UA9U3cos25KahgMITh/+4dsWDMOOacpHaNZdKnxZxeL0o9VmuGm
DmYKw9hDgw/qfXqcg703PgZ6g+fGPo+oj/PoLsG7b9JV3WVzacHwxsKoTIt4
Ujwe1GEORug8s+Knw/z2Nr9TbZYpVGubu9y+F7cRpUvudXne2Yu1dRg1IHRw
XMnv/u3BFwbmxWM8UZcq+l2m/GRikqlFb4L3asft9ZW/Y2It5Zz6Rb6RFsDx
p5AEHjyBXsvSxl2Rq8fVsJIRBm2TwmqrklcOF6qCywapaMOd0Wq+KFQay787
n30RqswyqeZGL3uSLAfVwtGWgOd88NfP6H2KkkkViy18wwpga7AAQQp0klsB
S0jeHUva0QpRWVYpGnorUPfkgl+nfl6D5Yi40IjZrfrnGxheojKhsmO+GBPK
lnNCRxIsHpMvf9lvzHL5/obO+Gmoi1Iy2Au1Upg0bqCYgJEooiFJEPyzndsp
Poq1FOHiTxR0t7Le48N9dCpQdW7thq6+mKPwFvy5J6ha45pSG16wIYEMgh3Z
Oh+U8geChyzedVQC7qqjtQK3jlEm5p47XpLvEhzsu1KAK9ubmZyjBdhpxIeA
kelOmsy/ZOC80VwayG/sJAKFePUzYUpekN6HTx7i6YeFzCXkX7Jom85XhxyF
1eCFVMTFrpaBVOCd8AqHoJXvkUT3C2ASU8iGRsaEghtTeqW+V5Vzr3UoKaro
rplDfWzkG9huJY2aTYx2I+5vqb95ODeKaKU2S63nR60F7aid0Lxi+e9JAN8Y
LcpeBQsF4sfqsub9CJHFHwfh5bAqSTfVB2fDPltaxHrPj0qN8p6klY6Fw7fW
05X4pd20SaoDvOgY6mqsNrQfasw1NJ9jDhxAJM+Lsr3JuKTDfE+Hc8a7qm9p
KopGFh5lbY0XWE4GmbXlybh0gWsqtjxU/IMhB1bbCuwwFrX9pkewiQBz1TEs
7sTG/Vd+WLQouEJZBGqKY/8uPBSj6ex4h5Z3JTLx1mKZJX6G2SPmKKBuh6V0
A4HC0oReIrmJlDZtS7AFi5rjnqN/6lJXiM+Xjg8IUrfqaGo/CWjKPdKhVK/M
B4NSTfV6HajOp6yQ+DEXyzky/1BtTJaPdPmIHYz1ZK8pusmb4NYy5urtbZdk
yQoQZ4WCXcga0xQRGspBsUMR1GtVXG7XrHkXeZ0sb1TbMKvMGF+82ihDCj5d
VQ8olV6GQSXxWQ4jKHx9RW3VJACubEE342uT8YUuigONNoKwtKludHRzLcrU
GUn3Bl8L2MR3edh5sjUzBUhvTwBav/q167sLgqJExZpxr1k3bsR5D6EPeixi
JqgYpnB/ht8eq1Q/p5/gJ+mSc43UVLuGXuhrfM65DDedyejuU1y49ToYg00K
XnRrYz4qFLlqSL5Neg91SBysh0geXhNUu674maUp31YfpDBT14YcKNAcB7zY
JWB/OKC8Yg97qXH3nFQ0ubXldR1udjQWjriVTQcQejDShmUJfXq9zv7B1J4Y
T4dKLBT/albipzev+PqLLRuKoIb0jsKrh0O4dRTWAI4wo7RlGijJ3A3BFun8
GXAYd5hz2HCMMkk8SAEv8bl9vrtgWPC++xdwMF06S5/q232ogx7p+hX7x1sh
WIXsu9xcR/Yz8GKiEzfHYyYLDIQtk2QXW87TmrSwzAIRe9C1ESvCnmkwEoi9
SFo28ldwsJkrNQ/CAWScPs0JBXPqR0IdJgp0IhEDBHaPudammTHbqT875rNE
mHlkyAxMKIWgry3hoT+FUR4qaIlwazT4Ceh5ur4S9aIYbnHeA8XFGe16vkEW
V1Ko66qXEcBfb5VQjTJJCRbWuvlqP0A0W2gAtbLjKbnmUUyp7G3EBomY80GV
uncwB40hD3dCNrhQht4RrT8ya7xKa7gTU3J12hochjs60mPcjHTNTVihilGa
QNvbK3AjUiFsMaE/eMP3+7VrUUjEUSomr4RKw1ZQ6v0z0Zr6Kq0Czuh5E4hp
EdKfmQ4zSla9xHKVon9JkmTNB7n1eKu6lA/pKegSxvlyfsTBjg15W46xpzZx
SIdu0x6+L5nYU6QSt3OUHGyvs87iBMPFOhE97Kr6S+JotLnv2q91R1y5/ajy
4RQVox0PT2twTj78SOU0T+v0blRW4LMj/H9o4lHVh2wSAp7yCRrQytr8y6jw
Vzxb75MvXy/5RpyZviC10cTOrsc4Dp7FMuymanrWuOtoDk/s5GX0Jz6iz0nr
h08EzbcpAHA/jBfIBXjccDF0tBZjSXih2YTfzOg+bDvscF3iHIHxDuytHaLu
yuCX200wh2IC5hYIEQQoHDIT9Sns2HEAJeLJHWgSzPY5t++FhjlhTG6pFPBb
HPV3EhNuwXntS062VfBIloXmV08PLdNhqaUyKIq0ckH+R9+dUsMuTWxbmF7b
XKlRPChkmmiaZwsz3qbQee3gZfsgTfxf4ko/iUFVRimZfoNzLNG4BTdmyN+w
YwMoRaJTO2ELTmR0XDcdOZ4EoYsTlEnvirMGOqnGJlvSVRy4Y838fnOw+xs7
hRahBnS9YCeotdilr2sAw9KJFKHg/k0RKwr764gOU0Jzp5+Mkwsgh3Z/BN98
YcJui0YPRVZuevQFXeH0c887DzSXEOKdHf6Le+zAi99zQfHx6CdmwrS4J/Rn
tKLdE9EtpZC2FCmiWYvirI9/v0s331ZbFS8VKMdHmd42xXBRSvzvN+xH5Ho5
bjswdn3p9XdmLu9YBqsIvO9VvFzzaXhtXW1IqTO+RAGpMKo+W45xTyLestUO
gZZ5nWyw9xp5oUCrPp0hCl/tYrxe0SpSMi07drJWpD7MAABiAE3SRhF0Wcy5
qqnwtNB9z6qZOImkIs6OLoEbmL3YoVmlZmP1m4KCckM32IbW9VYJIR7/t2Tj
rFaSPe3A5ONnY3y/M/Bwi5s1hyuhZBgEkpC7faOEvN5w+4BFF64vf3uYRMbE
+uLDgo62A/zQG5XYEuQY10fjAzsM/itKJ8nwd0H5eaP+e7OJcXcUwaEBZk60
I0KL+kTacpXPx5ylTzCIOsIGBKE3E0qi8+pl32CiT3uQXb59H0WZVOfnQRwo
N1Usn5UpFuXiGs9HSMQDuEutbtx+0njWcCXicaQJFP3ktg4Rh6eY6bYDuNqH
hWtsw2O48augVIakM5bPQ2oRIAYlYap31kH86nxBThuAW73A12C+TgRhs3XR
fAKWaUQQTzqwMdQKVITaeDCKwIg9lsi1KHCVjlE6EAEjucoJXnmtDO01k7SX
b/FweKkcw2v7UfooWoDyFaEoA2pn82qNfAJWI/Vk/Z9x1U4eTgBXbcJ/blpP
/vEcN8eAlEsCJkzPZg1R147GUAy/g0V5l6j2XBc33RzPan7mVIms53hKnj2k
2FHhQTbwBbDCAubTLD3xhAedU4ImNJDJI4q/8Q0pWTCJg2jhDRO1ZzANQ1G8
B/ciQgI/UtHUgvbpwPQwkFt7IhvoDQwKEObIG5ZnJdWF3CUD/iaR9CISEdAb
LVNTTtwW6sCLrbmdblqdoxIAjsZj68iXWgZEdFbo2ffJBREBST/QAddnoPMv
R2cv+wh8tnMx9JxJ7HlzDUkG2UpM/GTo6YqaLWe2y0+Pq8pnzYRdWdGSPHHR
x++GIZ1bujcesCjCBACkonUf9EDqC9z4e1miPLD4wV902m5Y41ctLUpg48bN
flLVAbrskZBpvoxK7VmSr2Uye1v+hjPgE/VBvjfXQO7dtYRHgNsuQAkwJ34b
5cHqDFyVxCE/AX4IxioZDOgM9MgwEL1hIOSbgmWyMtdKf2toTgmUqpll5s0Q
HY+7uUHWhDFBpSm1CGvgNrSlD7TYSoT81CqdCybTEwuR0mujyrB6XRXopmgn
GJNQz5wpWeVYV2IKfaHmKAkN2URWAk2GrJPsDf8r10NsEVdTb8ljvdQXZDTa
u87slSTU1Y/rMOmaxoV8M8lBvlWQZj4pSHplGQqJhc/n8uZzz0e0Cf++jIUJ
JuC+qwLT9TK4VhgN57tf3eUvpgmuj9Xrz4BG1/dyB/tGmVMYcubyA4fVsv2g
RhCuZkkMbFXll40z4xovweAKzmCpnS21Rk2T/+mRd4aGBQp4P5mMs57Y0nHm
EjpcuSlHSQckmc/w/C0/O4AxweQHWgw4ldc6PjGA9COOL80jMCNdCdOtfpu2
SslL+tUJ83fYdbnW5zysut+uRzjvKSn67Kp1W6+U9sxz6bXRUTrsqE+t2gb0
w5ukC0aDJ0a1zWVEyIXyoDFQiQAdnFuGzOSUlZyXPhW1Wk9Sj96cR54F9xwR
6FYrP1LM5SftFRFEdpQnTk03C3rrjrerilPrmQcUXxcnK/gtFU9plJHyocmU
V0CL/tLMerxh42yzLguqQaN2cJdiF8u2Mcu7SwWBcR9IDMUfI7qLFJTWr/ML
J4gzEXAHIf24uxESKoNKzSbEznb62lugcXhWcKrv2BiG11SUw+JKywFC8iAA
DVC+iVGf9Pl89GTguQ7LSOfj6qP+nu3kIZGSkvNOPFndLK7V+MI/dvsCF4MP
DKzxUwnds6iber9Rpd7bTrUlTco5Wbs8RI1P+XVwfTzn0uXDGSO4kuxsEnF9
I3bcdLh9IPCc84mfqKNoXx7z0ytCnXr3WRNqXGLwdkkFnf4j9r86QFwbPAol
U0KQxou6Rgl7tZax1cF8FvQGvl/0dt9rdC3eUGHILJFxuqM+wsWteJI3pAsS
kycIaCOeOZTRFkRcCl1s0tAIJtBYFmlwCXz1pbCjGe9vhAt4U1gImUGaGt2d
MWWvpTlZCvpBHWCwSjVLS5XWr5eTeh7kRSvC/DB/0qZQ6FShTeQCJg+WH3N3
roou0g0k7qUTq4kl+YHadXf68hpt/db4mm2kbBrMWt68KA3zI8XVnv8As2fi
24/oulqcsCxO7fLcV3hYJDeH5aIhpHPlaMMCwm+1839l0WPEbbST7UVKBtyi
+75BoVGD6zoigZYIT0bIpbcGQozidpn3TCnz1Dn/HG4+2T3Umx+GpMT7A7Kz
MP9iDYfVN0ap84gme4Sa2o9K3wvTYi+3PWtyOyGDmFuRQdVcrrn3sHYv5eYk
kJHjupd0xqtWDxJdRsPGcu1ng7IY6cWCPiVfqeP/lxjH3T26ttM+D3xAK96d
wAfZT107Wut4Y5Zq856mNzM6ajNEZfyVSqkTkZ0WzjdGq8tpfrUWg3ogCJC+
26WFraT5PH9Su32GqzFfg9n7ZeBsE8viPLp6VyioaJ4F0SRWKnkKbtbEx8Ne
+hUGOITEgbyEHRCqFKZa6p+ucy6+nWehON9Wr6Y1v45oPXUmBXV7EAiZ9gf5
6RXbT6rDtMQJ7oU7Bhb6xqr+ugHsVRyoF8nL+P8nRwHqXZaFzZYe1cYMoz21
7ESqxDMseuI3fPKf2RRaCrXIAj/7R2NoTwUp3xUGv7MGJjr8AsGCRl+Ik39C
GCXfIRWeJsP9oRPPu+tg8zrPBAp3is1T3TXw1KCPKYeEKZ4CizHzof+HfKYi
U1RTu9SC1+l7xl8rr80RuJctc3ykE3DIo8mAzGKcJ8A67wIootr5Nq7/VKLu
9IWfMKVPQmFvwZOUXsN77deBnkVlrrihi1WiACLby1AYgO9ZMsiRsD3X3K/R
5rmAMvYlWlLqqaZuUVC0vPtXFB8HGvJNv8i0QBjYcrlPwhGL/qBrGQvFVrgE
NWG69VHpL/YQirQuJpslrxrgMTArdTnD7pb6Y5Uytnbci3zWGNo01pDdgA69
ot6nOiQ5NMgkXGziEMpoCQN8EDtHtPDVkhmMji9vQUnT2lQk/AJb9MOkGNqS
YZ2wHo1wjIPkWbqaA+0ZTXCW0EZl9N6QpJVLsNKPcXIgq07KypUGVFHaCdrm
dm3e32wyWf9mkCAFgV8jy+PNjMgJYexIgm1opZ7K0Hg0E6K3vcAVU86SCpZU
i/wGyG6I5LH0zlTxfsbCIRnLvYdryEPiBq/hZgE7tVcz4wGX9PD5SNoh1KpA
MOhn5BSLqP03Prxu4vgtn/jiq7ObejYacMkUN6nKz+AAU9KUxgjOq+wcy/Sc
YXpV7KbSQ71HacMB3ScoEnkOn1lLtHuRyYmYvmCiN4YCpYCKIqNIKmdE+6Kd
rfJWPw7adaN7Bg+WMGjcvFlI1uKlVSjGkspo8Dw5+0tuta8atPDxHHFdhR8Z
segNOhVSjMdycZ9kodoc16WvclqdB1PCEcM+9FWAOpHirk4LEF0qI+q2lrma
B9fWrdJD/UR5IPa9tKVglcl8s4YG6Hz7sJvWseBIbRF8eSZhEFhAJNunSa1o
KU0ABJK0XY+Ndt90tllj1r8kXG7V4ndHdcmY1DRytVAPwLB0Wqum/GkiuJAW
LDkdW7wUgHTIejFijjoOspmwxt3oprJdIt3kviBp+B4kYkupiv5v5jdC1kQo
iUs46TPJszD+r9LR02sraC2EJdW8/Yizd+hJRJrlqooFA850WEJELVV9tvVw
MP3sBndkQRngAzR1O7VbeLuhM95JxhhTN4H8OjlC/V6NZtUr4NsuR+TcOxAn
7/N02EreeLERPEDyMF26bW3kO7Mtvw8a1+U/a0RoNImjdE4oa+YzUXhAMObW
5lpwNltWuthzkBdy8pihgISIIoYiK9Ov0y/iHasFfHH61t3rU2TksbZOe3NF
GKulWmwkjBp69L+whRQiXY9wU/DOCJzhA6JTFmNM8rl3hFmLgIIp1pNlCi8T
8ulBocKNIa25WeVIIDIgGfmt1EYmcFNjJJhcXDf6NjQYji6VzqDLucWTPq8k
uigtGuk9qXwjK/zQME7Hp0hFIy9vwqVr2MzRCMi8hamzKdVGK+0DiT+3/CyC
+NUrjwHW/NeV8Ix/NPr4UhD+lWUXs9UVDlGDPN8Gtz3EQxafiH2PyKT1WppX
KZFF1SOQLDDeHfCEGDqk6o4kXAbqXptWO6LUuxHLFYzS226po0K7pE8K96w4
DkHBCAVdE+CNK6wBFSnVuMurb+6kIimzmHajGo3rvi318Kn/uUSb7+3StZAe
poP++WE1SdPLI93ohifYIE4eK5JpJn2CeyBlhi6P3zsi1lH4AujsCqDef7ta
lcB39V08VITmv67uXjCTB84VCU6C3vjuSoU1vTEi5a7cH263jUs48KIV1cJA
s6ZIInAb9jE9GQ4DSO76ffX2wypwLPulSFQ5GSTF7ItOpIj7iqER1+rl5WHm
Zbd8x0pkRSNAdUT07QQIqI100UmCTDKfwcrH6a6EdKvNpEliMk6IzEOdwNT6
dV5zuC9IbvAvLJlxOhSw0a1627dl3JkdJMDj16237wbSKQvkzjKG1Vc7M363
QROUb25/u5fJ2G9kFRV4HBrwaZgvbBwhCJ+Dsc2dRvBi+sPZherSyj5RDsZ/
OIIgyk1yqv9dDy+Jq38IQTyuo57qx2dVYlM6vhbJAp4qA77xDZ8vFUT2XWME
A2rUkomyjZT2LRfjpeT2fju+syJiA4DnhYaPsoo1PI9RDMQaGQO24+w9L+zb
9Lwc6IGBt5dSJW9kCK9C3FFT4FWJGHVW5yhhGH3rB5o2AKx7dvke+sHQXHdX
wrX4cwG/TwOslLIkxCcVnph7r5bhAQfd8tai6hy3zXNmrDK6oUY/97bd6a+w
VZtVa/7iBy8lN7GoJAQOiust4NcIV+6pVmQ0ybIOKak3lJATo4nHH4M3/85L
WZe7Hk6H4RCm+FtNsnfWdYo0Quz2L2a9o7e4IixoD5COb3Mq4oPyNE6sIE7j
6e3jLfUfQGzDcN3bZ84ycIdgN4oIxSP/pY4nfNJ6v0RoEeKjhuD/VGJHcBvo
pb9L5drMDFuIB4GwsgYTMP9PjbrV7k2V56i/ZMguluMwanmm1dWIr+vXXE6t
PYB8ulC9VrU0LPRxqSShFHoIS/4CJ85jJ/RDBM1GS52X4xOBroORyfWd8XiP
z5bYfl/hrw4ep51pdK6h5Z6mrT1J7hAm78g/DE9kwhXr1zBWPKrN5IB/ssA+
5VFfLMpdvCKVkshzxa8LIVxPZpX4eW/QilI8NPxQkQHCCnRfWPIbbOPRCoY6
AL1v51UozH54G1fL4cC8qKaP/iYfO1f+4wGOqRq0Prpbw895KvWfufEIbHJl
A+O687kIvXDSbm0LaHNiLV0aUHlOF2BuXr7hJaZy79b0nJsrk7gZoJpC9K1P
0eRuF0GRJlylApU5lMnQzMKPOaLpUfDtbvw81RiMUfZVEsqPSrxLKxNY+DHq
3ZdkSx4zylFe/dG+mIze+DmYSHO0wa0q5LUkPDJ6A5vtEVpINWKOeNTU/MiN
OFN+ZAb1EVAxopGhyUQ7Y3pLyYy/urnPRV0lp4PoeQa6GF3yxqKon2QPzYRG
97Uj+VwTJQKQIUD0ghc+GgNDfDX31QZcBBwPLyurPlXG802Y53ltMZe0vx7H
45QuRR1J6bYk9jX2lahJ/2oZtLOuMcOTWmudxDN+kx2fJISztqAQ5Ro0ABQ8
vMkhCqO9VB/AT9V/gpuZ5qy2sAweXRYWG6DIoqmGKt24hxMh7CK4MgfVFu92
wtrIScvMQvQZtZSopyCEIyVnGWk1gO5BGzJgEp6OX47XX4Pf2rdkHKDg5gaX
QSZ6cXMcLBbWW9UKMjLieteL2g9KYcB4AREhWJzrn5/iiYgsSGx6WtjjOTev
qx90zqt5Qw6VVFVDEOb5/ghCmY5r0v29S3Dzy8nw4gT6/RDSeRU7S114ozw1
7MkTD0RWwE/Kcve0qidUgtyqVnAe4e/bZNa6s6uDgsihV5HZMwhOizsqOHG4
VjxPm0zBCoV+O8cBEm9VtJIBPtFuJWK9Cnqx0mLY9W9Z5jEn1aBXIJdUoRJ9
0Pi8zN+Vf7K7jlSmhPVoxtwTySTQBmFxw9akX1Nel3JGyvMmcTDLrLGAGagL
w1WagdkaPc8SsIMGO7VqU1k0JlDj8wrwI3Wk2vz9/512Q7cFAXjvz5d9Tvxh
EFpo/ZKqXADPOW6aQLwusmmTrrA45Uxljk4tt80y/p6wywIlM5QXt3hiwcBH
zB+IQKA9uFzteKgsOckAGG2jqrHCvTbYqOGWTZK8nUbuo2OjvxifDbUXJFvr
85ClIMv89gsRx1C49LekC+n7fZM0o2ZRWoJAeKYGhM2r/WAKsr4mC17WMhKI
dx8gOimg8Gihf16xQN0Jwwc90MAoi88UCsMh8s6RpiP0V09iw8otaWOx43a4
Y1H30iqMO9yp2k6kxsSLx9Cz+o+EN0dXB9H3gxUS9lnuEJMM2cJGs7p1BEM8
kx5r4b8PuqA70ioRL5jA+b4jQTie6xxvPniJxoUG59Fu46zsgiZr2Qz+I0Tk
8YWTgjzcCFA6XndXdyt49WaYLlnBpv2GrRWMoXlCW8Bzrdjesp1cY3IK5f2M
4Y9o5XjNOaSJ1AdgzGwOZQ2UBMXS7Bq1gLjLuvFb6CAoJQpwrk7pr4xy36Ig
2u/xswIcVPASW34BvqAPoL2jJJdKmZ6Qjw8EiF1A+JdQ65B/l9V4Uz36S1nt
ciZ8cSOc4II9g8QkS9A57tsVMnqFE9D6coxDsPVRc0+/9PbA918zboF2CA/E
Ny/pC11rqdwV+Xq5R22oM3nfy2b4erNxcOznvZ1mayrS2iRuqEBngeCjr56/
VTU314miyu+r+NzzhecWrYQGRitZk6MpaCijGLCxGX8VOSZpx3dJp3Ygj/lL
ak54UbfT6egeV2QK9U6FhEef3zu2ktkcKqASrDm3wJ5aCqInyCiepOFZDjyW
Dn1+oneM0jXbgzF7tVqkqMA8Q1P2+snnuJ0bupiFTBmbYp0Nc/O1LlNXPcZb
veuVj+PXf/T+eq/cln1REUq5IRTQmjpNxDP4nhUfmR4B6X80LDDYhLTTRT2h
EtL6kKFFj6vLKu09Plt+y+ydwyDPO0qQ1g0XwFSzx81yF7UJ3ucBXjZJhqyJ
ezMn4HltLx5HjwrmJwkYes8L/yM+PP07GK7DkM38sp/UkUGu/hihCoaje7Ct
7SFXlCuH3Ubx3WMA+cKFxgesL9NGj3TmHgGm2Kwb9AGG7hHnj36c2SUbL1yB
UEWkkVyRySSvPKwAil6F2tBakYuv+pQ2Xavg8i2t/WXjSxwCW71NqSAWq7Bv
8mllIZnsd8wQc5/nhIeTkpd6+vyxsAMtcp2eRcRbV8JjLI4wE/BcACqGBBeo
23K3oscWMCjdC3GBVG22gkJXnWbtIl03qmayjMtan15OnpUDEKYfsfahgNem
F31FZzqiQMmbprxRScpJicnBghjtCZl+0IpXSubKegddJrS6PkMnJa3PtlR3
Sn2do7tcvrCf65a6HWr5qGDGN3p8fMKghcdlmkASIJUCi/CeixQ+eb876QxW
Gslz44Wm5W2wwd3nM7szowUpeDhPN93h/ouud2nIkMFFBPKbPoZudjlIFnS5
in9PA7n5gkNfKwzi/C2HEWprPQub50EjWa/ZIs0MRz/fdOj/akrJ6wmrWHcu
ggZzNSRVOPez7TyTIe9K3ewWz53a6xQNm8ZRHOcUVl9pXgpWWy88rtZw783z
tWOrefI8vUDgoc26RHn4fH09W2/UVBRnS13ZGJtArSCN26bTA8AgMdiLJ+U+
z99JeI2YfVX/CbDM4bftwNLiRuDT9K+Zy4w51FsZvcK3SzF8raYajbCPIAtM
gCzn4KCLLa/yvBCHKHI8Cm/8tv0lWW4FhIvmGlfATNqSiM9sGsNxXLstB27e
oZQVTxosMXosrvUnrH8I9s9MX8Fk8LBRgpCXHylAZ0zh1OvsoSI4LRoshX8k
HPVZrk2Cq3iu/wq5M77nij19kc7UT7TMdvVE7c8hSawXaZslStxscvL3QM+v
o5lp6yt16lzLLnlK2N+y6rBIdrgb7Q1agifgGM/Hsuwr8TYGmh4JOwOhH7aB
ZCc54PgzrcPWs9RtFq5s0/AeuIYQGeoiXQkhTasHd9xTJoXSvwTjubKon+K0
gm/soQiE4Nwnc+HeU090bgqsqvNxTC/cMnrzRZ7aYR2e7TtB10vrJbqlUfGU
6RQYtfeSHSzO83ywRkTAcTG9J+vN7BIhVfq0Y3AcpLfIrjbdqGZK9jq9Nr5u
2t96zOxb5EI+JKazv8+T8wUyGQz/jM4axVbGoRx0wPe8jDvrTYOHtnT0Popf
1NROkeNdCWfaClVjIGuzYuJaNi1Vxr4hk/5xWKEqBR0O5ajX89tdr+AKFTwH
g6IO4BZCQNewwpS6ZQFRxe2Z98rpmW7hy3IRcw38JyQQVFF5Kz/PJOh+roOz
mQLazR1sw1PFsHRJpUpmA1/XsSb54cJk7IAIVoF7nGnTyFGHhXxT6sObYM86
kmQEOdBvuhrYJbSV7bzCV9EDv2bk01dVNsQDg4vMiuLvQr3e0oSg9j4eiEL9
TGPn7PrxSpo/NPZwlZWcU3CEw2wLZS12fGdnatuhRud5JftZ7fCJ5HE8/RYA
6UJO2HdyU/eg/jk4lldh6ZkmiFHWBw5qszZAL19QKH8bMsG5uWez/A3tc9lE
lBYFdT6i5WHo7sBxhpOkc0/+oumbhCY+OZOMrO8LaRGRmu/KvpxH2ZYN99nU
k+mJGh/zbC/Gryk7UMU2W8UTOr93EHHvS8Ybii4U0R4cehRUplBzo71yyzvI
V4wuwcxo6zDT23TM/3YpRrb5mtvBrqi/xautfo2DyT9tEQOuTSzprisdUdKc
rgfk7fk01D63Pm9REkqOonxdRcZg0mmAuCa+pm/9sd84NPvhycWVa96FbhPD
1XVP4p0MueC8Pz0Yklwd0OabN8eAS6IsucO4oEe1IMiAOAejt9C4i4A/qqY8
ZGpdCHO8dHo3DDhx9ziFGM4DGeNNfE1/yF0a0GaNcWFpaEOZw1uqn1aLxwlh
rLKhD9/j/ng5/7pUhwCU74Sjm9RRiYUl6nuQgYHu3a66AL7ryxT6cWN++2bS
Gyeooa+4ygC7X+XRl2w/izXTX5A/8+bWbDmOA6pPgumdp8PoWqTvwOef15ha
FCgAfSnu5gkcstufkKQhS5gLSwFYq6B7JgeyADXt1+MrO+nskkb4D/deFLSV
uB+qewM4ZUvZle3rP6npwsEjuU8iHTT0X0h5jgQmkeOn/fbUFMUu65NOgYwp
TTK28F1fpdd5ALpds0W9W913qRs47juKSgBikHpjhfHFEpmNMU6MnZvbQ7bn
4sv7iqXLNFR13RoyP2lyCQ2xSetc7iMtTYm0qKxow5P0U4yPYdbnp21jSamN
B1JHpLkCovdHOoXO2vkXe7IaUCOstqST6jNm3N7db0fM4TqEYD+oRaGOwEqB
93Z/uQH11SmO77vkw4hYTJDZg7pOWhkisR9WMPzMfVPWjG7hMi5bItXjDRtZ
BVm7UIPO6M69PGqEeU70XaQxpA8a8/GKAyl7HQGZ7SRwSzL154IeYnRtBBqH
zuryP+tpxEUeUddl4wZSmiyrx0VdSiDZ8mEIyFOpJxUMRJMLkBdXQ8gLy/DG
UjsyS8stvsGf9XFEWeM1nm9miJuhuTc+a9dLFUPOGjBIuHyhg7p04aw5i/EP
reChv9HkPP7wEf1v3rcWO8OdTsD1MJSZUU4tFDqgJvXyApXTfr/Xr7nW7JOs
0Ji2StvUXslYJXpkCht8SGrCiVG2xDvuta0IysMvoqJX9CbdYi4gEjJYiKVe
k3j2w5eL5Uv+gerLxg76t1157Q22+CcBKKPwt/k9Q9g6A3WzpZu7hDBFo1CA
CD8gHxWDj7Jxbft2ky3vso1O3aRzMJ3C7ZxRu3jLadsGQBoqNdTscw1w3FWs
vvCoM6zyqhdEw/yzVMGxdAZh/Rr6BR1bqswHmkq4fXvuuA8iEzfC2mzWqYI3
fZ72rFTuEnKZviPcoXaGmILndGwsrj2/bZzAX42Y5HWCTY7SdLggK63UEQMK
osg1hSggmSVDudsyFAutRfKwxvHDqQsXTxSojmo4f8tqyc2Aewl/VnOJBN0Z
VoZUBe/7fmAZGSVbl/faPMe3VpEGuRRyD1ntHkpIqyUyt/1CLl6DW1PPuh75
Jor9hHMZqGXxz2EYauyx4nCW+2Vu30j7S1y5wIYuBe4uZbmwItBsjW5r360W
CFvijb9U5pot0SRM+2PsqfI7pYJiK9KDobKfgkEJqPQU4hDnJ8iZ/Ua5dj/y
BLB3P0z6q3b7/cmcRrQiog2LQoAC/SXJ+6NA4PKpGKOZmDISMSFCnv8HTGh4
eOtjhCsLNrvZKwgWJTNbpw7kEe6NJFBAIzUuIbiETlL4zJNLt+m1sDTKKwX8
uzI5d+biWU8yzWgN3yD6XRBaFwcMOZreHAcxh/Kbai8zZnykVoucAJUAkdRQ
Z5PjrMBxqMVuWstPbEhLYJBc0spGxZUmztdFpFzJ6s8TBwZmA90ujxxzmLaB
7M199azL/R3MeiL0b0VIO+tins+Zr2OBCKNQfcNbO+E3rsBpr5XuPesPpmtr
0Cv8z5ZEAnyax3hu92u2ZKs0hjumqf1ZCXoq37Yxm/PbpPNzAeiUnZ+zgaAY
NpLAySpCLEJnH+CBoj6y8oEEPQdSm5Hk9oe8CgI4k5J3mJApBgYBYdy5jQlX
/ONcRGYtfsxy4FuM5BjkzUdkJn9lD8/O8fguNV56IzJL22YNESGaGr0v/VLI
vsGBYsyvwCiZeFu2tpVU/U8SJLhJT1jzcWDQMEZ5LWK8gJhkargIfmJL2mMq
0pQD64AESJ3t6GHiHTkiv9a2Y4/D97cBXMJOhncE/6J6vh8QT0JTJ2hmUtbC
rI1EUCuNlUEPE0uSPpaJrkcPQubkGKKkjilhd13koZRuIuzk9pOdDAVvrzJM
hl3gDdo2Z33fuK8sUj+t5kRBbrs13cL5ki8gQD/UL9tROtdELaAoT2Upe99A
oBtBKYL9gNrejI5XNKFS3m+FvXBnkcWSk9/tfjF+mBkhTIMPh4FGXjLzxk0f
IlSexy55Ko5KBX/dsFKqcK4eai+eqGAtF3eJ6F1pjHLJIwZSbTb8rpnMymZz
04f3m/sAvmxFm8Bv73VOyP3mPWqIX7/MX9zKkj7ojaWQdvOskgSVquC/BxRN
picrU8ZKesVabPtNjpjLyWgyUWOsUYTMBorQ/VMiqRhB459VRmJER/U8VA+W
A1d/g3rfxa1eAhj7jqlpz9oe4vKUoYcMcpREq2Ig+zHmMiRGKC3jFnZZ86NK
S1u1q4YXstuRmIU36leoE/uyGTVklQrH+5TCvmG6RZCw/eyF+IPmu0GKRTfk
KrOm296QrG4EQ1Uh5+DPOe1AFnKTKjsG1HYOCRM7dK2+QL4jT3XpJuD3K7Qe
h3tYurd9sZDGmtYEu+yRovsPXMRTv/TuHbI/RvEQksehIJl2JqQH+dhQUXtr
Ywc0nJ+NLRSYPChdt+ZOje/D6PqAcSkr5jPuSJU/4pqT2eguQsMM4rq7I2Qh
BwatJRey3jMkJgDxWzHaYWRtXhr2cCrr3vWf3h7Ugi5H+2TRWIC+8tLvf+uK
9wqXFa0kXTQYkXN14VSgMrQH3ZI8exJAsCwHm/kIMWLeyC+CiailfYw28JuH
QMqhGObRzlbMtQfpv55ldkork2qkT2mx3cbs+BWcq1YTdnnIQX8etncxdNeG
9e7KiT5g4EPd4wt9bz8QehcKf8uFkLsWy7Ke+xYTMggqnY5rcT9NVZb6fvwC
bJO2kYotkrLm33IE2FQfSUzLuuHMVWhtgjzCPx5ZCENSVD2ZDE/IFoDO0p4R
5IroTW99sESBowT99fm2KZyaqxkiSGCaLFQQ6mpLhWfvqmaSp3W5MT2DiDPM
sySYCKX1mtIQLt0GGOx0cDRXWlWc0SnBFDsWAMhJa4wqyQ2W2JPyJU/pUk44
MyHfTH+Nv5yqiCFdDuXrNlFwof5AnTHiu9YtSoo1jKS8De7vx5ESTOwnZ7QV
BWt2eYr2yu8wqFr1fM43tud0rnJ2CLkYZzhl+hYuyXXmAAik3wJbWAxWSP9h
hvENP+NWXvwKz3sDKtfLs0PIyV5DehaC0bsUxudM3VNzn3aHz2Mj7U4B/C6s
SGBv0at9cWwh+qbggvmCaI5DfYN2xVypq/hYpqX2wMsE5wYPRFkHI2V6DjN+
1lPN+G7YzfcL57Sm0YVSiRxuJZQ71rL02gvXQrBVGscnFVVSe8McX5pwDTb/
0ZqMsP7prijvSzEUgkpBuaOB5HlaIgqdK5Rarr8NU7f8wB2y06bveoLEhcoB
D0zWllFro6pOo0GWI53/dKBZ5fND52gR0ZmMQQVW+g7QlUICXIvonjHpEXu3
rfwQ4i+BADLuMT9L8uXAnrD1nv1iAsLMzAJzSS71OVvTbDwlSua4o9k4eoeG
LGrSKS/9HwyhW6OfBKdQFVqvkk9u2lrsrYJFoyvvFz0lENDVAPGalZaphRIs
/sqENLbLd8GlVjgptja/4rBAXShskWoCDXYj8rzftKBjeGOEFib2X7dKj0J3
SuVOJTQEvd1EsZdj+MwyULqONlIJjBpk2p+Ghi9G6ZgrSeCOQT/FOmWEPjBe
cB1COffkTW6/blnQ7QNWbOJ4ZIKjx8DOhfmpWaXvUj1m28NLzpqFwWLg71pZ
wKcj4/cq8O1QL49xIUnzucKlKdE+9sswXXPCTj3G6SHr0YXoGIslGgLqG1Pm
p8aM8bTlswBmYzfMTXxGj9HyonMs+dek1a0e8QWzaf6dtaCf1dRXeoAgq5+q
UvHHA0ovZPenQRXVIi9BZurLrDNlWFsD74bonU1VT56vWPsyh+kyjJ8DOxie
i9Tdwo7sODMuL5DvTwB/wsApR1phaz+Z+acYQ+W+FPAMMQnLEajD+B+D85wr
R/F2IqipYcddMvtjRy7FtS1eZ8Z3peT8zGTRgpPcU0sV0uQ2v6dWqEtQeiMY
MlQQkYjVrCS54hcnmPWJjOtuwQDdvc4SBozV1GlYEXyZB+QMCNIJYNZD3GCz
ZQKS9y+WHAyWrzgGTXErjV5s4NehCh2W/FhG7KLdzqtGjqK4EM6hsgh99Tq4
mGWiWtSJms8xOJ3UqXoYjddXV6uRt5oqzLKcD3HiJhhgvBGfRw0Cj6r0XyXk
RS8Cd+EWeK0g5/HI/m6rNRhPIaAh3tlUYz/0RxpONs4CVn6qBBiyC7maq3ZK
xzShH3lYUXbwe3mmHhS/i7Zm36lnFUfrMmtGrgxXKsdBAtV0/0UOkOuQMZSe
HV5frpw7bIqbZvLMlL7b8+ugZRAfCnockflb79oVuvEDYIpsIL5u5OlwHEEw
n7iUSBSBKVUqZgxX5WbAuxno9HBIZRgjzqkrTlzdpPG4aRMsFdQTfQPMTdYD
NeYx99N9dOwAXTfF0tPFY/qJLsuaaDiDJ3flpkDOf9k0NVgMsnuUXreHk/CX
xOYae3aABsu3NbIuQ3Bj4rbHwqhEQDT8YEgPWzo8PE9DlzqTvmFFbkm+uzci
n9z5tgkMOoO6JiTr2GlOPEVRUQYxEr3kOPTL/Ly1H0EzHQpPFjawY6Sq9OPI
WHujhvBAtcO0Ufaj4u6lAZfXpjWFV7kzT5Nh7+IiPOCmXiJKsSf29pI9NDKc
XnUW6VCQio3ywmDLGEELDoVWl1N9izWh6lhdmV/CaP+luxpkHG8was3iOhlg
9hJvToY2i9b4EpFXIdMYLyv4v+rKJ2A+K000OQOQFDaiO0hfRxX0job+mL9P
5VI3RHjgbbBQf6VrXQGkhGyqWo0NQSnPYyC2XGlbDqtsDCaoRZLvEzaVaRVp
6XT3Lv3TM6hXj4vfX4IJg+KwjAMH5ITi2c2D4ic6c7VlV9d9PKPnaa17LA/z
jk8G3Tbwr47Z4oSmkOeTnbGfE0/3TBS+0Qyoplw70M4Sxe2hFcClcB/D4OWb
VYoL8+r7ZYmSbi0yl4nT3BnexKN7gZHuH9nfEZUlrrA/i8NKsiZJKviJjgxe
MkSZxZpu9EYeRbV812ohEqmdWRbOv/20D5g78Pb0mt+6WKlkwMq6Xbr8yf+p
kmJTFD2aJd81EJH3M/w+xnttRARRXpp5ZIPTgCKgDvTbHfI4H++QQs1s1OVg
erpmi5mPUNLkbmhSyvCmSN3M6SYTack+2D8SsQi6Sai7FJ/LojYdM2p86KBl
o3rzpBLjEPDXfpqBWDWi3FOGXAhGsOcR8cSl5iMNm1bTfju+yl85bnmBt1Oa
kVeiGhB8HCzKrsFoo4ZFYy7GYZNSVzXNpXzt9ZhFE8aPaa0GV/iiC+bgr+a6
QsG1Rsm/wO+UVHg0mOhkNeXdBDfbYAKJGe+k0cZMeuVCyCK3oYh/Gk4zp3Jw
UbLqAzUhPDkmvxjN52yKACgJufPsuZ1cxn+hAMTXMc/veFxpRMiW+pN/tL9u
LZoCJYA3pLwwV086glNgOiA/+RjZ3afDhzsD7aZ0riuO+EWbJvqKX4ShhhvD
YQPFdcynxPDZKb7wixYYYChORjPIZ0OgNiObwo/fdBq14fXHjjOdPqLPrys6
XgTBGGvWEMj3gKRhXueGmhATfDcviopCIL3q2KHr30ytBcS/q1JFUnf3/ByZ
/bsDOgxqYWYGRZqLs1UlCHiKVy348LyqAJRipAb0H44IVBGKfEIPcbR+v617
wEQov0Kw3xZ+sQrTg08DC+FqDrYi1IsezbJhYX0w7TW4KsBJYcMar9mOigIg
Qm/DEOKxVFU6S2MIy3MhV24mSLDwquXbqfLc3fRzHwEbGJuXS60FULM/jO0v
k3yr7mvW9IXgJty7JNWvaVro3sMdejhOIa+BZqSeAyKUir/ki8GCmqOhyKU9
M/aB2z7yyR971+L41aAv69q/8CItWhBpIuJ2yXQh5MTKmquMJbtHMhjONFhm
6yQdtIDSzPkxmDijW7v1D72hWD1j/ZcOTvbJzT06I1BbqVtRf+TU8JenBAOs
/lZFKI2hmLtb6ws2mEr3nwIXqu9jlf99DyKbViZuwciqdpR2JL2UTxjPikuB
P4YuqS1PCmR6pPbXrqzveE1v9bsk6Tr5XPLrIc1ZYk3bKcs6hvdmYSXpTYNK
lBq4WxbP0CFcSoevt30xpOEY6ZqD7D4aqSoIfLtmSNGy0MqSH2IJne3ktRNi
t4sb/mRivYKMOlyID8ewNZAvnUqaIMBSv3siEvITMPIyMRTJ4ayMcJJMAviN
oCE3tAuNlc1foi3b80+RjMY9MFcVe9GmTd7SUIRcuq/Ofj6FG/YFuJOUIaGi
jm8RJ8/bezW5qITpSrT4o5/lHT0b5RXXdOAXX0IN/dG2eJ/MtIRmhqnCpZb4
cO1bNIlhcy3eawryTaGROMzO6YE+aXsvEIDSEVweE/5lNHXfe/g0q6ceBOQr
3Cgl5Oo4T1WEOOsQyRk6aul+PpVy53FJzttQjKUR5Rt7dTvFVipovmNptoNu
enXyJ5USI/xtX2nx6Qc4LrXW6afMAcLfUcKJQRTpL7uVA/ybyIVpMqXWT+GV
a/F8NZWdKEO0UE8sSclkGMoETXP7sYXC3Cp0U9sLSiXmo5u3K4NUprc6w7Ds
sURToyW5Dh41ieTwqnV7gR1WGizOpCPwoAJfKer5mMEf3So3ebyIeSz+fRYu
8IOzIYosILCd472EkEQ0RkIh5yAWZJ1a146eJRexpTPN7JXSu/NGCpcy3kuL
Vtg0vse/iHp0DguLq0HBOgTOfjZl+mZzDg6RY9TP420SL/39r/0qAPKMhrlE
4GxSE6/p2nqmGD6IxLHTMdu8DcReNrho2/FFKZoJM+uGRcIq1Hl25jV5uOPe
wouuya/IBLgkzOy2pYdkcBOnS5CPodE+MVyPBJVgb2Xq3RUq5zyohG/29wMw
WmeILnch2eMFe/TZK8TrFAS7qhYUw6iJ4jmTqW6Wci/chIEfrlQa3zFAltJD
BXzyb0C3AcISn3Y8IWaJw78kRN4Wyc2gI+Afldj/JEL8JxYX8OenBWm9s9QN
soBQNX+3qmLE/ZBVH3tbdQwTdDFlJa/54vpgecxJkT6bD/FBK2l7PBUGQHLI
wSmaLw/1Z+1I9NFctBdcVt2vAQW/L6YNg+BTNKIdDTK6PphaigQIOluBJa3I
UfTkmAmnENYhLo1BQQo+8uHJLXkGhVauCXUXAlD8LmETP6gaWRSK9yWFYo9X
9bO2Nc6P/XL2rLiieA5ZpJzmHjw3lhvytvS19erxdFVpvCl1CbD4UiPKqvSb
MevSa3KDU2/YwnGiaXbhRTiu9NnSUXvVUkG9NK3lLUZw8120C8V3yR4zoGQR
tOwYKJB+6c6WUjyZY1eBRR8iVZ2pN4AKjhfN9x0nTt766QGVk/XCckmARF6f
YuNf1inVs1Ohfur7/zGTZYH4IgxOKFoBgJYctOVOJG9XKKpDlFpAU4LvLqdH
ba5g6fCKuNu8wZPS5YmWLqWY2afgPTvIReR9hC4OBb0AMRnO3Js6e+dYDf0K
Rg6pVBs5ib7/03Hk+lhvE27SMhQ/5WEaWyDlgYPT0P8MpVDZr76RVVxfZrwx
RisXfONkTta1yDdA2MqmEMnftt3YxDbB8hPL9uycEuV3ak6Js/tNUO89vrbr
/EG0ruMftk1TQM4wisQkow+WqZgz92Hs1KxIf97pzCnSRcNaQamedjLxIbPu
lVUbvY+X3tmVFNc0No/Hak8WFC2DcxurGX3zJ9ORBqfnm3h+g/EQp1WZBMgv
h8iUUuFBGgDFhpO+x0sKSd7f0Xrujwox2P5mR05g4Q5pz0DK/SnjJrURNnIV
MSWZ+pS0JB+UKmvq+o4u7MH9evaXyuxP7DZeeTdQEEmPnT8IqCxpjxMIsooQ
XeAoT0jT5gVZ8XZtBgToNsfhjfc82VxVxVo6biZ3P525gtjp2RFLAM9yjlCG
8AWPJbYf3iCQnVf5aEfXoIs8PwLmmx4bsCIgrmYgckY6seY0lZctYUqVFtIg
36VGrBrWjWKTjwIYrl+yEqZQtv4AzqqE/uy7JG35t53wnpLrqi6LFlkvd7F+
MTp0c4Ew2vTEkvYqeS3ni/UdO8ELUkNyvwR0xr99OWBkazf00YKNgMOvPr1h
RyituQo8ZU+nGAvTM25NmuAzYhenK7G7nqPvdAS+06SRLTZv7gg2VSidBXS3
H3R09FFJHZk3UyQ5OeWGt+qBY9E9sU0MNY8swwI46mB22QvrBREZxRK+NWu1
CehZutgSS7PJLOlkDRBkM96vvSCK3qEACH0+jRNMRIKOtAreurIwDeHxl8H7
t0l1fuBW0dFkwY8rzeFmfZseDpv/Ycu1Qf76BH3sm0DlOCZIznqjGCm84566
FQK0K0hHNxJoqaqntawP8X4NwpIFTE+Ay0Th+qC+xZ9e/j+QbIENR+TDwVCp
zd1w5VKHIv9sYxz+HFoZYSHBBauaW3TSRD+EyRzeWIKZuTlzscLIiuSsCnfD
woDxHGoOQenWEvYXDahJVdeq4hdKvWSMR+Y9WZX+BOZlNX2c1R5V9fgWc4ja
maTDLgtIuKLUc+MKvYpZC+DWRyfFs0gMspmjgLaxKFK6N3NSSj42Ry1bXgxb
2Esrja5wg6ytIBtXrWJ5bPjFSUcZJuHG3WL+rAtBtG79YRNCr3wVJsffT11a
UY0tWOmnHdy1boozWQWNwLIIF6VbplaPLsNGEt479gp9Mf0Lg9HQprFWwY1p
Ew7g26ZihYIcsQ+HuGKYck7TZWBURRxYJjqTz5HDySRmglug4OfKp1/yHVLL
kxSt1w1yXzfsReZWdSAyBvjlVBy4EkOrdlU1Qy9EB5PjNCp/II6L8J/E+uj5
zHpegRWK2l+bPXXZmshGXvnuEPgX0ATvatc2V8EY6Qxpj6Ne31EJcv+N3TGE
J+0oWGRl6DiCHPiPZ7oXSxP3ZEpmzAtOQK6BCwNNyeiAWm2yyFvNWBcKRqbb
y6Akooy6kvx0GKBqSLJl7o+SDIITxZgJEyhK2xdh9SwKkt9RJLpb34PQUoXp
cUTpU6cfrWGFcGVCuXRYU79m+bzSQIbk+Al6xbL2TkQ6+nDspUdii2irzbqM
l3QpxB7eL5DfAg6E+vRT6vgkpFsiHR3rcPpA4eI/oACe1jyFkbgA1RBUScH7
lxwj9iyHd8fzsSBWJLDZ7CDOq1mApNLZcymZhb8OPFzMEEDDF4dQAv3DN8g0
XzotXRcbvMFaLEPUnFo8y+MW5py7Y9suTtBBe6iIn3i7xF4KUj1O4ssjXSsQ
cxJNBBFIYsdhr0w6+N9hEgnLaLmIuCzzZsfej5v+i3CSy5Ycz+y+2yRVIqSB
7P+UTI60S56FPpVio0wcTGUgTbmJ2t4XaIfLlDklc48zVV5ROqOUN7k27aQV
CquFdLDL9z0AF9kKmj+9u+J2LggfJnZt0csi2JKRwKX+Rb7/q7e8rG3S70H/
93mmKktoVFVis4Vj6itFDCrBwri5yz0a80v6buMJRoC1Vn0e/9T/6Q1WZP63
ZZFBn3eyVE7hrXeogMlnUHmmmiPYYr7Pcv6lGxbyp09RUveELl149hEIvk6x
Zhi3B89QfmL8VJo5GsS1MTOQKwDwLIUBnpVBS+EFHcLWkDcIKlD2yHzJjAf5
Goqgg9sZojcbuCxR7GgDCs1wTYEvUK8LCUiNdgzMQQlmBf1AmyaL7TNJMmfF
EKWjqZwT96J/uUaBGwbGuwxCvuVPlSJi9XR6tEsvwfYlkOeVGw+qu2XXg0im
m6rk7sjOH2wQOaaSD7EKXH6UeO9O+hwHW4rmB+KL4k8aTEv1958kbjotRX1B
kwL00AmFbrNDoNCt38jhYLKRcOQkvHY7fOQd+Kw393iogpPRADy2dgKfOlP9
K2gcrpIk+U0T+evosrJxAJjq0aWXLPrh6+oPJ/qWO5xsk0HV4Dui9tIAoZs3
nJRfFfeU+RacFGhf2R9JYdi7UBMcT++CGPHg0+1Fhw9U2fkkiNqjjnc/DStM
17/icSBU2n+ytqJrd5TY3iIggS9PbdNkbfGAMxAU+BMVKAuAZ1TNfbrSS8+t
irYa6W6ageBbMDoxsD8SiZZ+KWkBP3/svvU0RaS2FvW22sNo2Int5cX/GxYv
Ac65aMIoxwG8Nyhu2FG/7Da/q6uAEy+bUDSrZnqOkFa9NmCjxt7bn6U0wysB
pPaVWvA49fOePAdfrIeJJIu1TJN8F+0o9ELyt26DgbNd3ljhR5HyJdyGceM9
YPrZ5Tdp+Le4MOCpc2ZUEMZFzFul2bmS+FylkQqsgfOWVuidj/8yWsTZY9OV
PowFkeENh4pVmIP8x2Po3ERilEcOSJl8VfqBgUY8rCnmb5yqhWwtW8oDgPXm
fO9WWxdZOktIOPWRlc7Kxzkw6Pbky5CnSIlbq3e99lQenzUYUPQEs7p7E5yZ
AilBb6Qvm44pCFhvkF1BKoQ0m/X8jFObiH+0NStXKV9woy6jI2AjHMf6BRK6
QvO7mieK3ezIFTPQGkj86R07dD3BvOlmmGvAvbY8ETgefPDcJj4JCDy4OOFT
gJD+Id0svYCZyrwQuYPC7ImB/kNQj/PgFNJom0VsPvpTQOA8ATJqBFomg76F
1niDQ7WBRMDEudlx+40oPWOPSfvehJzsEfUc9YJJI88wBBJSix89+qfMuhX+
HQaiQfEdQYviXP4lBtf0+pEPdm5H48PCPANndqqzVH38BBFUQQ31/V880Kr3
5bn17//yeSG+SLMY2HY67jARiq5BMGKl7xLCmhXTZMCgmqhyaj5gD2ZX+goP
KL+KiqQF6RunkeVHuYOsLMI8Kf0bkEJ7m1dC47EIUXmdlJcOi2VwtojFfg8j
KkkXm7m6M2iemSCrxSsk1A75KEnXJpQhO1GcnkRzDH1x06f4YVPfPO7WuOHq
/h26bBmtnlY7FmMl8XWysZyAKbuawsvBVqFFJOo7luN00NYeNI4bHYYQ3ePm
s5rlBgNaP8JqZlaoy1Unm/yeM0jCqM2KaOWIzbe5VNxcv8/vvK2CH5MajcTf
STa6z8LbzyZZwmcINCrn34MwHTdx1ByXz/+I4zvlL72Uhkmdw8Mk01XSBTaV
I8ky8ARv1QW7W3iH+F26jV+6ysKXmBhvC4rT4YK0Rvk5Ltrtc8anqZf8klUB
z8am7+b1pdfADRAnt1Jf5TFbB638gBvZ1Mddx4oLgpxVY6vmQNzB+FRCEt6B
ujIP7iWSf7GpMJZyFuvtSuOguYhef9yvWr1EzD2jqBsW09nCUWzcd7tC5KtZ
XiWHLjSemIqPraSwrpLkZgxEoREvnLESObAgfbjvfw1avSwV8EOuehSKpxzD
ukwuatCBXVgQknn5JRl9+VENy7mhTI6w4rtuflm4Boknfj9va3pbrWbZ7byD
V9V9X+28wR/Hun9lxiRGIwZRhKunxmYHCmtW0X6yiV+9P/htxEY+WPxy7xhg
m4A0W15RwoqJSaYKv9YVOildnJvcpU/uTIKqOMT0Yy16cp2PSty8W7jTj17G
YVldKe9BlcuPareeOnpPLlABimQWfOjpoObuJRX85YdWnPKr2Mr95OdAo/9m
88zyYgqElYD17p0/aoeIwSzBmKf/HaMwd5xWWjIqEOCLN6b3Ub6HZt3Wzww5
Z4J4wiw+7xypVE7QwLgh5hfScvORJEQWgKGe50zO524kFT7eIrMV9YWkVemd
TKcTjNWkoPLyiOVerPOrgL4+X6++LbrBuITLc2a5gkJ0Jx6pOeUNOVk/92n1
ZdV8+VlMaT+JBb8h6kOOXarGwbSLoDbFIAGrfbcelq8OI/coefMvbNmPZed7
hkKyxcDdB4mXICALVZQ45i8deQw8zY0wThri5PiV4yKdwxVFhQDWyUwEcwiM
AuGf3aFfl3dm4vcJW6kSHW114YrZ3Nh2vLUzTflejBujYfRPh9lWSrOSfPS3
HzhI7nmJFhXn3hknyIOrDVpJIlIp49ZflKmBUW8I/60F0lTodiKuN49L19DB
rei1ExtjDc7qQ/FEIJH5lb0PP3u1HuF/6qo8XqvMg54x4ERgsKJ0sq0SG30P
hCkFAO/eaio7vdTevFLU3LrjmuSZlVuyveD4YTVD7owCEB9pu9v1ZcQGHcJW
qRcAC50FnJ3mwU7w5aC4rnIO73AnPxjQXE4bo+Wo9q3fHiCcwoyG+IcP8z21
H+KRWzR/QygPEDFZskSO3hPr4VIYovnAPSCEctEOWmj34AQJk91ItQs6u7lI
IobTkNcpKW/5UMB+QiFu6cwOy5vUkBP047zNUFckEi0HO+awpMqIwUhuMESG
03ujeepasIxy2Jqgfyd1xyTKfErv9EeE7YTd+c8dTbzxzmc1wFSPIqg2lAWi
WZNBAisv1VFLFXOosSuHXtQQDAK/KlfePUtFlkO0SR+9geimBtuB76J7qbHZ
GgWL9AMCq+ZiJFdt2/uS2nbbsolLNSPYUQn3j36f4Jft8JU1wsz7xfNCLA9s
vx1h+cJ+SuxvTYpqeA7HBmRGy5lYskvKR2IR6yCg0QEB5dbENmpDhnvywzAt
2zYLsGKGnXlhVS0lN/wiSvWD3YfCbzXbejbMBjsz5WSyAILeD/ThTjljrNjG
9L+/lTHPaWJMmgfBhSUsatz5GDk0OqbUxYW4A9DzOkdsF7FHlSl9XHZzfUw1
S8s4ZZt5Ol6y/T9pPpXUMX45vuT//A9HxW7eFft9cMD+WuE+lpYIUHLCzbak
cQMeFZhBVstlsdhcOg4q0P7Fbc7O/wG3zyBrosqk08DNineC8rkwqwdmLdC6
PFv/N6APXphte9tQzFeGI429noE9DX3PAO0IwootI3z/gknG7fXc0B7PvSmT
WUcEvy90dybVmyu+URL7y88gIZo5kNB561kO6yj0XVtqF3fc/wnOTeW7rrRK
rOEMXULTJEodE0ww5cdZ3pImOuAQy0DCDs+WVC33XPuNhMrnJkOdpCz4xYff
Fl95rWB7DkSoUj9kKsu7BtMustqttIimz7qJkGwW0JWWUiqO3N1w7WMTyIOc
RRYo2E4+tljO/onXpBjeIt5bUt6p/yIx/mx121Z9xt755qnVF4UBvII2uNkE
i0BqJzbxZZnY5y0CGg34w+ym2wsFBL9Gu1hSEUmoH45xq6TG8rH7KBbJFIJ0
Hg5cpsHLM/8y+fQ8UBxJMjU6uaeINe05A71MAV29jKenQi9WWDLlo2Ho4BRP
buoSPdJJBmLiu7HxFMCXoTgbpeYyajUBRuWVTjogWhhMOH7aOHib7YjJ8acI
LLUPurZoSycpy9Zib6Hu5r253EF4NLiVM/r5tgar1MlEukKzSvDTW7djmxBT
XAh7OgJvb6lGlIZhmnTNpZkhnB65Sv1YJef5qUHqPTug2qRVlpFDePyX921O
KVECZ+/pqMViMqGap+RsYCrov3k64SSxl3p/OKQ71R7etAZm9LbWyWSbHwA+
7CceRoq27cE8vSkNfiuCDhu1mkKX0gRHaBE0sDYEPawYO/hEuVy+i28KGQpm
m9AqJ6GMAmhqOjdfeHzXKQusIE6ElLn7rjloWfkY+XiZLmX+PKmwWbrvPjrU
FBo4NTUs/TbdqNxtY/b5UtyD0NRxUhSX7CLi7+Xr8zlDy2kXLPEFgpX7b+n2
LRj1iLeMDKzYHN1HnU6bWQXyvlr9yh5umhsHpyOwKNRsu7w9GwcGUy+RtdD4
qxGoffnAnkpJP41htH4QerPQ+C4dJQRuPZX9k3l+4t3SqLkOlACOpHLNpZ4u
ydnDb1KRrbsRFIdSIiyItIFvV400bL0cKF1y/n+uZgeonuB3XcCkPJZ7+u+n
9oM8rTggbswHq67ULB+LueGwqRd5t5agYAeOCMWG62g0CXUYHSUwMkqgLV18
kj36fPrE3dja/sM/h8Dj4mG6WjaBc5T2CaKkCciN2vRvPBotvVIZ6Wmi/gRU
hJekphBmd/+VjFdMz/lLlYAvsMF2u+8Cy/eOljksAxFzK6AcOZSbwcTgL5YB
NJ5V/IACYszzqVMsGfvnOeV5nbAuRm32Etx88NM2ZprCTeNtiP0Cr8vAqMZv
qtInEbue5TG9Udd7Eqzl9pcpfCeo+rnLQ/YqvG4H2FUBvcjdflYF8eAW/cH/
iuEUZP2R5m32fNJc7fxWkvzgwGJuH5/o22fhOzfLTE1V6LT1vBI54ApRj30K
rWamqV8JHw0/lj/FttTt8wlfbMOGmWgJExMmeR4ml9JY6/iMr+EkO8wxA31a
nuapJI/YxHMyV1RHxYvf08DFYOo+Kwukx3t5iiNa90ETrtBd9q8S5ErMhIQF
gxVe2K/K5gMYi0cxSqNTa3o5YgQ2QTkQNL+nv4zkgvbRxSsW4CymvoyATjmE
mQcYHtRrH0NjiB0lu3VkTQOJ20/8rfEcl+Jm3If/aSmrSKIDOxJvMBDn6MHI
qnblA0oj2xOJ3eJs0LgS3hM78UnKPu4Q9FtGhbx2Pj8yf46u39uZs1yAo1vo
ND8DK4V4AJYxIJpBVgJNLK6xth6UqzouoNEXghBUjT9Dm9tSZn+5SgKmHmTg
mxLiM3oQd+wTVHkLUGWZpbaZRwQn2RYZ3E4tY3PE3++5x+R1D4J2nhxXwIG6
AErVrfjemYirrr8Uk5oeC+gbZ3iVTaoCoA5yB3ID8q2iaT5HGYN00KoCF+Cd
uLOH0wCPaH02cVjWn7O/kF51zZUYE1iD9K4t36HoFIZecVCAXL0IDcesaEIa
Sghg7jLYoCgnGvW7r9skqIzRFoq4uR5IsIosSuJXRTe4e62JWzTZXzrhiIP0
m4+p2tG3uPpvNYQkESBsz5lYScnV8nI7QBH3FoLQ7PEiAr/5Ln5/BBh5zGKV
bYoc776RuyEnkQXM45AsCKzP0JaWM17gaKx4n8paApEJ5GQVqHT6+Vtu9haR
HhJMHxw/uMIsXsWgfJcCXlr+ek8cbadcPVU+OT+jq6gGYarQSij/zTC+9zW1
UcFfYYN6NlT8Ym9tL9CY1Wy+V8hKnuobBhsCfmPaxuls0aUtRqjxVtfb+trw
yUQjgt7aSv8eHejAwLZlQitFtZ6xRNQFhPS7ffWoz6FJN2+EXJk/uxQYd3Xc
+bawUHNnjL7LBFdkc4mZMZWF5K0pHw4FYv6AdG9uu/J1+QmRBWqo+HtvW/NI
hzr4Le3TF6wOm4+UBjw5j8uy35k1VaRXGWVE5SFSsX8DpuhaMNdGmWP9bDV8
AT3zUAzb/hXJLX/HlXz4zqT9Q+ddCAEN5Fc/IwK0uYq1l8ww8S3AdvLWJ8Kd
pg6QEIkHFgjQbO9/qn0RJiWZ5MLUecsWEHUd/pKY5XetPO15NC/UJpripk3w
Ecmt9I7PK3XKJNIeHQpP96edHH9umSn62H5fmAr1EtaKm29b5nZxz2GBcgIA
822HYOMkoVABVpLPnlkA2rI0LrUdcviKPJWLSR7nulHMHI5Ki+97EDaRHW4d
e0tWPTbsCvcFFTf6i87H1N+FmRv9VNunGxW0c2q7JuqyU99O8Ali0GpRUqXp
nY+ptjsNO2e6eeVSJ9bLbqoUfz72k+fpbDH0WGpoFabjDO2kYyyvN+C6qxYG
c2yo0WrozLblJmBAxL5J7ripECazk/1AsQsk+rlSlv0dVbJlzC2fpvqrJc6+
85pgdDdTvLTH7suhtx46lFtXO5y9dDfFQKAARnbvFJloOq6eavGUfKH3Ptgx
DOausZ519a/ZZy4H9RKp5v7dqhdRqj63o27rLizCCnDASUR83XpPFf8cJFuy
vcsUQxhyKt75kOsFEpatBT/5P4aNFPDVYQg13TnYXL/WmR0Vn4m0cSEarhZ6
ojQW1UIcdxxYXoqMJQpNNYKntpVDLqe8mMlV5CfauVNUFGMCl5tszfmilThM
h+9kjKk+YDPof4rNRQxYrrF7RJI2ql5iazBJChWsWyfH8E53XQ36n06hdAyi
nZjSPUdpZQYq70263CwuTNdU07MhPMq+e550Eaodl53rJVin2e4Zyz86nk1A
2DtYMZwpXaZXVKPIYY2BqLPb6N1H4VBjyY9UlAxMABtSpnrbrENMnO6MOXRA
GqgXZytDQ+IVQfZf5xTWSQWhdiWGQz0C6j78L/mteW9ODPZ6f/nUiKRX3sYD
hoHYwyw2bX0W+Hm65kju9aD0lRZ8TQNLE3UFjTascLHeFxW0blhXOPnR6gJz
pyvxd3aztgIw2Mr0c71m0nqjg4LFfjQlPvnv/xTKH5Z5nuTi+T6NWhgg44dD
c1oIwv+6fm058n2Sas3NM3AdrOxHDhOeCrygYJz14GHSTS7d+yY6bm4Hedkk
BRd9ELjuQa5J6RKJNcZTB8YqZDjnrceodIxrK/WnQkcZ+1Z71pwbEJJEHSf1
7GQ7O8Xc1q2+8cHXtAFFAkiT4opijfNO3CwPKPK1Rc52lX9/3ovb2dYQa6iv
n+hMKKHF7NulPOLCHchGjGx2DuFL/bR2bBnw5f8f7r7i9ICFTPCNb0CKPHKZ
FJh15ZBYRnSBpfbxRZ5GX0VBRAiDv/oe5Reb1E7CzwwL0LGIqMzJ7EggZfmJ
qT3tgARIRoH/XcgwZtXVsYLeeu6XMssU3u42K47lYE1CQQPpTNkI7Gmov4j8
8SLoGJSHexlxb26K/A0ebKbTOmR6iJKfNTy8J/aqbND0elusjTM8uQlwytzl
rDznWti74+9eAk2DW8WTpDyNm7U2bj45keUgoZSPUj4k9ZdRk1Qq+2XfvecE
WuHroP6q+uBNb3jaBMsZ8gLT5SUBATpCuSjypM19dJzlfZWkLNxHnhe/SXo7
w+DbE91ppKdyZ6z2IUtLiEwUyN2Fdt1dpzVeDDdebMAkhtLiL6H0RTQHM2+O
khCtyv3XiDIdw7TTJfSaskZD7xdcGtP8qDvJfadzSpPvgpRCaYIKQ82l6mgb
esE8G1NAVuVab5vTqDrVVtiWtG/I9Qu8c68Q5T03IdoR8wtDJ3FzuYON35rK
962Pf6Ej+lJM0u8bVPJ5pHP1Q2+wGRWf+a5NMSzDzZ/eWzGrlPtOcEcQa9In
P7IiINYDxLnEx42UGQl/IqXBFD+JU5iFLHdlqgCCzuxvPpi3MuvgYtEBKPhT
g/in3umAUay/zvfrSOX/EBBFNgMBDtcMVpGLR4jC6qAesuLclsV66lb1Ee7H
a8xSmOIS3Bw6ESAtC++b8Z9soEuPqiyMLCHrEfQkyCFDiTw15zEMeCTCMO94
/C5RDRrp5BISGFboHXdHfg7yfrXQHcTL72Sgd0chakLGgQ2LTwHy9xDcSrwZ
+Ub3iLorHG/XyK798fEcP4j0vaDDZssUbrEs2NEK4Dfc2+wAIrVaFyXgyQVi
1GgWjkc4HwGuGIp5hZOyHiCUJ2qMjeQslC3FBJj0818z5OxgWB66EOyKFT/2
BLOgcxyjCddzMNKs6t3+nb6Qzv+ltysuRQ6DaI7U7RLXIeRsUpy7HYCTuhfw
h5WHp4cOeANohVEPTjBTbOv62ujafhstZAkV4KXDseoFs30UANUCw3CKk0lg
FtsmFxMywgGCxhdDJKv0rYC8PQuxgVIsSOVkQrx0E554IbAU9E9r9jkjoW2B
bbKD8j0Ko9yw0/FExeMxK2M+q0kU4VjWdI9gY0rDF5Knp3aGaWpFYI9skEOB
vSWk112OSLKb4SfTPVAJxn14cyCeq8yJcD8cOAWn/Cr9VZhXkbrsqN9QEdvI
NGsLrSeZI931+tVK+0IvWILbsq4vrU2SFRfcpzJKFCY3kwDxrReqtxXaznwX
QlAFLiDJPSdzvtsxtsuEJroS/ayj0S0WK8k6m6CnZkPXckWUcMuSjInr0m4W
p8KffhEhsK15l84uNrU9u9Bgwx8hFgPPCN6OeiVwS3vCQbWt/7rZ8A11YTg6
rD6NXDlUhqxCWQr3r7Xn6eNuoKhCn/RYNkCmCYmGXDcqsWtQ/TB2/+slerab
wSE8M/uvm3m/yNylbX7aCMr3IqaE6Ec9MzF+TbfVJPoZQuoAAWoXnFBl1BLw
wc7O4JyLqwOQYhzDGDDzKF7g1ViGaWNq3KFDplWPM8Y4ExvKQY5eJaCFXP0o
qAn9v5ie3bITlKW1CO3iBwQfPSwJaA1vKVUsyU4KW986lhp2ccnPkB88Nj5C
WPB9TYoiCDAhKbbDd+pchZZ8VqzYX7BDtH3LBDPufIBQzJwXC8YaxHbZ83Rc
FVLn7OALjDC3DZu8hmUK88qNtXMIZda0Ur62arl167Nlikac/8qrbA6JP06z
E8TJZF/w5i5B6xoiS1mmXiKGs5CeDxRW9f5GEeg8fuqiMJq2lrAt36FeZBs8
c5WqsUsXEFeOYgwarqFCsxdB1OR/fJb4wR9Jcjte1HSSgsIvQCaRNeyZDTBi
UbtRH59FnlFzNd95CvJPRLJVvCPHIoX7pkhw/VyqyFGUl/y8bKDLCGtDv89d
B1dPSCnqW1yA1Cx95h3Ddq2hmJDuy+XehZ96N8545xqjik+yJLkS5pOs30Kz
Z6BZjcYw8Gvx/ouECQTVBSENpwkg2yLdrtTIBQRhXaRh6XreEpHFYIGzE84v
oTpdicg41S9+VMGXsNLnltP+dNrNVeVBIxvDMF9Vpsqz9aD6qibrfNfqW8XK
hVFd989Wrdn+Nb+IdW+rZseQljNStq7+28F3U5zUlOaGVxDuWkc8Rm8MDctm
srDjwqDbdlXMnqQfeQODNfqbDFjBBA3hmYE2dAPkpxFeeiyfRFfRhbBnTvb5
stKcNU9+pu6LcZWKN5ZwXGkKvfba8QuY8NwcqSGINawHiJ3LeS2Ko+pmOW0u
QQgxCPzKP0PDQcbErqNH59ahrEbqWbK7fo2HbYy285yQx7T70Iwz14g/MnNj
rbq3KeJqqsJLNnhm5klDMuQY6KFSu/dDw5Hj7/4n7U/vRZ8IHNog4D6QDIMD
GARL5qrgpz8wIiq0rvoZH7WXaF8eFI98fIuwJiBGqLix78qNuGzs1GR81iM0
qPjBQPc9ckxPzLOe/BC8gURx7NFpyuPS600XOhusQpp0Wreq99WHXk2g8POi
mKi4YBqa+HeqGz4L68ZwS+lDqX7sKxZU93N7l/Fn5/f9eSolYWW7YHxnjKfb
ErN/OTOgecoo4vNdJM5EHFYZKL5sboF7n2iKlrG8kLPEFUHviiRFwdmyNLyP
jCAzuZKOH+A3n2xQ5kxWyOo0U1IkMlRZtAam265zyVtqA3ompZpo7wHpTrvW
esXg0egwD4e1DoMakNgRlyeSeUranEeER3mEXkWx/vvWKXDUlnaDkNyxptcE
+Irx6jmi8JANbFlK1fFYh9WkvnN36xYaRspPT1H+Bc3SWDylcuhG4x3NHtha
4Ons/4gJaoxHCM4B5undWxG/YNhUoN0oKifWKdhnx2uYL0mMQ/ViLI4UUEdw
+97IOks8Q4XUxJEXuBEns7kfL58jFx/HKE131ZGsXrXmfZ0hoLlilhXoS32W
uREcGyJetEDc2ziK3Z0ogzQa0unD8YoXbeZSwiEHX7qA5cqTXh7KdzScFhfH
KzxF3Gr6kQQ7DFWPs8CO+hRGucagn8qgnyDe42Qs9BFerEoUUa9IuSlz4IAC
AHSrvMF99cH9pIocdZxT2NrYugHFKr2tAqnSMIzR89jNB3o/ymi8Bo+52A7e
ZFJMOuniEjC6j4Z1L7oeemXdsmNSLy2hOeCb8EElPwmDHIvS/0WNZi+YUCxf
F1uLQ4wrQQkcJA1TSI4bGJp9PqAsZvxg6iKD+SAEDlJWE773bLKy9pCR9Z63
J/uPSsJvpYybbc6utr++iIKSzryT6Ki2e97ao7XNApeNnlAye17aIyNMnzEs
A9U80GrbyUHxBfeeOqBkHrfz8ml+zOZAPzNLdQYgOFzV2os5UBrXk+qBxZAY
lZV5aU0n91HGkp3ExXAS1lhSTFzxJ0O6cHZgUBA8ETZ8g9lrkhC5+PMHwsMl
O4hL6BdKo4GRbLrcJkSCegErmW6TQ1F2otoYKZI8aHneBVnebL3to1kTeFEx
NOHPewyc5M4wZsOkr8eeds9cGyyPl5qvl0H1iE8ew2iZnY6iZw28Dyh5ezPU
Zvl9mAxISVOiDZz+GYKsiX48zkmb6VVB/mhqnQWSK68rJ9K74U1NdtkaPzUz
dUud7ic8S04I/9PyIS826aKucpgHkGPu7Hoah3KRqezxVEV48jYCygo2yveG
P3jJ1M5uN1f4ubUK7uxSfki0Ldeym3odckxeKSMC3wRHXFKwm4z7Lm03bb6E
tQld9fgA6RFaxzUMtn08KBL3paq7aUUTxij9YuxEwmD6GZ12/gIwkmGelPxb
MqqL0W+3jEl+pEg8hLmSBDXKn1aYz2u7sRgw7Fw0Cy6RTyvtsR90Oz4eJ97H
o+lJnUvCubiDWBU+3373Bpe5++K+qK5UCcrLwnwlLJJtC/5N9K6g0Vb6y6D8
fSE2J29u0tQr4dBfFYyQsXOqUzGJEdC+D0P5kNPkk3Wv1OSeESTsFciq5JR1
vveC8BcAM1nSNAVXo1pikh5u3O/mXc2FJUvJbYKyPvokr6fZc2gesy7AetDe
8wkSDz8Ywa+HMvb8j5Zun9WW2yXu2aEmKEgK/Qr/SddpDhT6017iVdbg9wx3
asc4CgUhNiK1gdriYVAV5r299+LCExLm6ncY8Cjp6+Y5fmRFjKwpDxUMw/+X
b/dStoDEQUkxIAuf8BCsKPanbq45xlIF1NiGBUNooppBCGmH6aa0i45AHTMG
ckfGKBGNDxMPsX8gSvDBOy4ZDTdkVdLC5gYwfs3P1K83q+BdqWw5opJkRIob
ZYJXnauxNX4F7iMiz95u2WAxSeMGCE3NfTkzqv0qfQOj4rMgVIHheqzpE/SI
R+kwaRMHuvXItKYTNyNBK0g4qmCGWSriBQqZpkemt1QwF3lgG3507TPMLWHL
e8KoUUjGomjG5Gc3kQUo3nt5u4IrrZS/g0Db0CmLcePzaq/dnnSpD6WzmkbF
D+kYlF6Zf+CdOVca+Q0259g01h/9hpXttOE1c8gCGMc3ezz88IzrjAbb3buJ
kH3ZJCHRr+EJWgt7b1gTS5eJDNRB7OMqeuUCzcfImno51CKnF0WxRQYr41bt
Fkmc/2ctW94Bg/Yke/8mG+dcTcPykuB6R2Gfgq3pt4zl35qSX627gPAVwe78
pQlZpr2YPIfKiuUSZo7GvB+FfNpZZ6ZXdB+D4jz7aaBezKP2JoOW4KJVn7Pb
7Gjt0S1VRy08oigEXlvgCGIe0vmEj9tgTF6DVs3BMjaBxVTFg3bxTy6QLFHx
E0OTW0yiStF8SCquyy7Je/F/MIhZoE4ztMJ7lx7p34CuvXlkUigfQRrecodo
XzH6LwjJzOIlA++76W5hJtbb0zgAGEVo38njA49Osm66kcZqzJWewDnc5XMz
TsQjIKgHqZ9HxtshZRYsoax7VQA4pxrMJ3jHYZkUe7xRZttG9CVsUEBimj/7
OZwmrmQvhMbdogn/TAG/PzQHNrxKjLuOI6ZEBTYJrLHVPWJPEYHRBvR9pGA5
EPrvaC3Lev94I3iC0jMyaR2FWQx1EuTmK/xaRl6GKBth4UvH1Fw1kCsIQZRF
DcS7KO8oQ/J/v1WUheGN9Qf6UHekffrhIwzuWETVCWmEb2nMpdLsJMqgA5FJ
yYXdX+88DYTGWZsviUe/lOCvy59TjA0ISoINY2/sDfYTRZRDkgQHw5OUcckZ
LAKmO9spzqNrUTbz2p5aGeBjZKaPD6F/BZw1QtFzvRW18Z7Q3SfmkUWa5hOL
kpEVN3vOq/mMMOvArIui+wBtHL1Od8fa/aChrjA+sumrLPKQ0aB87U9ISCUy
FJoUrITTU991JDMmyHRVnAnyMuMh2cBHBOcACUoRaZd06t7v5BOUXlkXBLC1
JoJm7NTP4X1mruzym47jUM7m4Ruv1P7NW3nPbHq6ar0EyTkbenpznJGoFCVK
i5rGhuy3+/ix7m98JWGCnyHMvmeWrWPEcmitW+9WsGfrg7lzDL1+GsyzrO3C
fglBFSt2nKb74oq9BCnx91BExAQQabcQJ68JVbRajqVOd16RALHwqKdxJb/n
24EcNMdAOEfOimcvsi3LZ+jdicRg6sgwirEEReHL/3/X2sJNj6BL93NEvCBv
6PqRx5KIR0VSCS+hS62uddP7rLwbC55LI6kG4N3ULB4aqXSahRWelVkHwTUD
fgE8xVUOSQapc6GYwTb4hHZwG+5heEXA4+aV0e7LnHkYtXUk1p9DaSsO43j7
jwD0ZawPwS2jrZujvRjQVRAJOM1jbAaw4YqWMAZH//+cT/GiPFfdhflgv9Y2
JAncl1jl5uKzjgs1o9ErXfj10WzvYJB78L81m/pDxjf1ifub3E8U/bFjdsr/
GGKM4dVeqtBziEmpk2ZDh9kGIgp1c3XimDqWW8lzmvsgnvJJtU6bh0+F+3eS
8VgpAEqbttM5QOsvuPcZ4D/KoKxWwPnaDlYidxyk4yIkPEBt7ndR6HeXQ1Qc
TJkVsiDlDb1WJLmpDIJTm9QqTU1JzBSmTRDdiplWPcTxmgEeGJtd8M5s80A4
jWm4Zf4DnY1YFlRdVVwwulW7G1Wwsq6vAJl+c1JeRltN2bZn8wsOydvxY0AO
fYRA+Gnn0QwrY5k2fLE23Ds+bewIaEPez5a0cIJ1tIjau90VwQzsg9ZOcNFv
4jdq8d08T/X36+yOIiV+eIwrdebEIyC7ZhWYbpkiUZ7eXhde+sWgvxplD2Vr
qJ9JfPctdr0zb/BSrRM6feCJsnengP93RdNHC3hyaQgebSlfru5mBjH4zcWH
+TIoWRXrKx5w7S/Q+MgKbqtzGYbs8hOKEuSskwViRPd7FElqxr7+5YA94ue0
zrygap7h76N86I81cIQ3+loZGn2Oq1frG0VLE3MIJ/35TJdC+MrqBreBxIya
xWMpkvVO1lu7jAGBr1gVLhhiSrNlcWpteOnGxB/luFkrcF7JG4L4VWW/Kp6K
R4wo5deXYIrof/27SlT+nh/FYdi4zfj6v13gGIGsPqeO72/96RK8NBqWATYg
aspVGBtkVGoDGvftgCPNipwgWfy6M9pfkjybCIVbf3xSY3GyXazDQ6elgQCY
FqdxmMVpozTq6Q71luV3kOLNwzpsvpyyzh6ejgWeGW4ooFsvk6zq/tUg3gBW
nVxmh13SfJKqxyAlWhlL9vDTPOF1qsIj37y7Fg1WmBbOyAsLTWmnreWue/Jz
h9MawxeGmhuw6CoMwAD3zJD0OQ9p71zlrrunCQPA3cGSG5Ig7zn1DeA0grO2
VcDW8/QU0pP7QK212O/nwDQei5oEqUDs7ufbxU8DveUt/Hli41a3CsXMUKl4
Cd95TQ7Gpy8rdozi7mm4KtDyJV7zghtN6+WzcC43V1CB5jLn1VEIbdvcUcdf
w88gk/4Ex93eY1EZU9poLZtUl/k45Hzuoty1jgP2gH0Z3D/ztLxAMtxICeM0
P23t+Tum43PsC9cqfEC7zNQqIwGw3wZdIGwqTrVyfmMKhj5eIWBuCLMowu52
c1dTiDgcZCY8tuB6WCCZb7i9I1/Ye5greDwOvXK7+sXsgP1rjaf9gDWPvF8j
Dhs20yu+r5gVpgSwXxR7zOnBSOv9BKFUzN+JbpCLTjPLKIwUEYCPbGQOVDsd
v1kcNT94BUdxsUrNKBFOXUgG4673jx8gNIZP9gH25Xzj4f4IwCfGvz/JAP/F
5XZ2rzbY+0chLKG7A77lJrw0YyaYwYI67lHC4rwU6+CtnUF1Igm8eplf1JOo
UOkhcUAeVzxaU8jMUB69tKuaCz447hA9vwUhhIMJLSuDtumwekgvjHI7FHmk
obnUvnVcA8+nPgtHKFWQp7jyZ7BFILgEnkBbmW8sLDjTQ5tx9zf8cD8drZ4q
AijL9YFBVvBuqsFb5oVYv+5LVqN5A0HdFmYD/7Qbwv6Mwan+ZtgWmAqHOg6n
4FwaZDcbbmVTs/lIUCDnArGdrq3rISZL6kvjA2SVOytlevoEn4Ukf8wzkET4
xqBCSxtfT4w3k6wZZ6A2ThywOUYcZAK9RD5lMC0+hxDD011huxzRLejT2n0a
C8TtDndyjyvMhkmYrBNw1wHCXGx8KI39OJ+5GcPBuftZXR6ek43ZpVCF7kKH
PSpjomMPn5teOzqU3T7RcRxpdDccM+m1K0JSi+5LjMxexZEbmUlH4TVm/QR0
eanOybx+YjPgIC3IBS+Ckb/SNHZtUkiZ7N3R0X9V22/7l1//5M2697uCJOrF
nFNj6LMNNrUws7YfPWy01qHd7pPat7uW+WjwEJQdhDRYxjaQzUD49lB1OwwR
TghAbKnW++5Wm3YBY3gLngVkobpNtZjsnEHKx9WcrEDGr6gNSYq1HaIw8A0J
r+4o440SIA4oUlcvg6AOezV8hNzyP1gTKzHNJ2QbC0FPTss/M7bhn5NXchjc
bHelKAY0w1TK3zmyfREcH2gMd41RCpRMSgXsoZwhPbiZBMFuA3YEAkYSnNT+
dFFdIwv8wPGIiWVCFSjxiMpBRbZBI8x6oQsrTMdvTbZpEkYDYfnIW6n6F8l8
cS4+BQo3wC27u/fpPIzze/5vNd4tWoqOu5ZwK9apvfO1VmsNHp39l0Iobbtx
/1uUbDXKzO3Qzje0VUf4jr/BPhq/+xVA//qGtXrjhbJ+IkblmOn1EWk8RinU
RZ92IRqFxSr8oSIKOohIAmhaqAp+33QjL6sYP2kSWqeUiY/2KCuDbVAu/Vjk
bD/yfhLuVXaSlu8KePXbqnh8jxvbeGfGxuC1yvrYuvwOxAMQQxX/QXcRKrz0
5UcTiBsyhRfjTzIaS/1IwD+huvYUXBkKSnTOUlEavaOQK8wfkO4l/6C0MdCr
GE5AYqvMSb7IjWfzWJDFpGxOekccXEmEsvKmYEjvanjupdFpTpNQKYsjphhc
ssanJPgo3/uAURi1YwZ+L/mNTa7HnBYoPwl6jTctW2MpJrqFlMziF5jH1S4+
fojlgclHiaMPxcHTQVZatufZrtZV2NWHsXLM42KrmZz9Tm/QvBUBaKrBy6d5
BneejTzBTQTqaHpQzxZZ0KssSIPJjC2P8FCvtomtHfblrQLhM2v7xlhEHTjO
4Lk+bk2EEWMDLBd9jcssL2ms1tmQhOXnRT+Wzw7zHN0TeDF9RaRZuqOvyxfh
dmHQdX60E9/KfCTMwAaTGXN4jkQIO9rSVDowm563ncbsC8KNN/Gfu6vbRlPy
eUJrFAzIeOutzmNf6vysjk3I6K/2n4qDKu7Ixy2pg987/A0AFdLuBLQDjK+H
KCwg8B6dSPlIHscTDIjsFWPlqfF2oUpHFDfRFWIB5SogGAroIcl3i2+rqsFn
p5lJl+URG5Cym8bxKd31G1fH1YpyKMEhSPRyBiM8Vd0HRuFxvZt0ylST2r1N
sHAEEN35si7xpfsnIdIxsRb9xSuYIDKhjrU+r44WgI7w5yIa2tEgXY3pk/91
pM84MMTD+BHq3Rvky/Lr2D+eYbQEc0ndXJ26L6vZnMcYKLkDwURwxAlYguKs
qcSH4t89FZh1A12cKgI7SRuYd3H751EuAjkqdFik5tHzcc/6broDNhxQ10Qu
lwzeSgzPziQESrJjgmQ3i7f2HErQBg6fkn3sil3lXp3ktuemMY/w0lQuVtDc
7pVM3uFZOEChorn3lz6eJSGZmCe1kWxPbzvXqoiREbuGSIhrMoLo/9BLGsHG
alwaWBJwsEy+Md6U6e3gawfrREzWJwE0b/j4GOKzOQy7uT6ScL1XO56QaTOF
GCUe/eKtXkBpqbtwRlADtYNVNNoOn5z98I62Xk1Vlj7qyk541VZfbmFEzbgJ
4dcrdFzZIcZ3aq0U130VfcWBqM9/CwwSDxWtJ9noKhkdjqbG3Z8jdGvaPv0/
kQcOltjw6WKC+5ZQ2VqxIyWnqpG0Ymi6NjlMGuWhf8RwxMXpja1iBRwPx0zC
2f13zVYf7ad2VtDmWUZB4pnNe+1xkMl9a6msGnOjr9mM1vbboUoufH5crYP7
AkqYcri9wNyPU2TREQ3dpyv7q9lWJ6lJ4NF3BNjeEYQgFBedp0Z/Ltr26lNQ
GLxzE4cXRdCYZB8Gj9SvF8CcKL8oCmwFRRhZIR0OXJbOxYCd5iET9CjgooXH
OPYdEnPMeF3foSWBJ/MpOmp7MefkzipZ086gZH9JhEnhdiffqF0y/mRBE7jf
8Zum1lA8nrUIJjUzahSmr7GaE5uGl9tIVz/TGmjbPjJq4oIP0h7+3n3IH6EL
dKDtXxjXaidLekY5O4/UhXVbc7X428SXcc4Rqk1ym1ux17xtOfcrBoDC7q9F
G70m287GlkVKcCRgd/kxoclsJ0RyWQXiEIUouv+awBlp9jGd1p8BjOP1Am/g
5YxtHSUD4ukmdTvowdoNa3jEsYAD2VchRZ+72ptLuBsVFp1IB5GvbGXs1RSh
OhUj2ft5PB/oE7w99xKw62fUCfbH6S6B233Mno14YHycreCiTgVkBEzx2N6j
L3KRJMkHhxK35L7gwhdY+Y8quPEg887Nb105clQJrRKKWOvBzpDjcQIm3fv6
076J1IwcWtIBvAMMWeq7z3A77WcYuKbYMdOqoNHGpjE62nM8x5EG2CIgI7UG
Qatdz8NBd0pAOdAv6oPC5g/gYqprXp17DqYjMFdSXOgHb8Rph3rjL1Exmfkg
LPkxE1SwfBj9EEiEaXQZVPUraQTMiYNx0jy8qaYb05RmrIhGVpT3IBR1J2YY
5DeSwPjBCmxJPfGQZ30xLuzhOFe1JLs3Awa6g1VelA1IC1fvotSVehx/AUUd
mw6fhfK1ojRwQTNcQ4QxlW/GJeEpYbFsEV0IdYKptv1PAfeURklLdGn+DZtQ
+B+k5UbLaCX8eOP4sdE1NBuWkiUANVReXrbzYm4pvnDt+aMWi1ryL5ccZpBP
Axwt0J9sLbjUpGMKRrvKdqge22xgVt9gwgoyu+deT48W3NI8h78yURNOQYEt
Sd6vtB3mgqq6wgN3r/thwBU/sXuMe6Wjj9n7ml398wVYQmHo49Nq/v3jlsfs
iAgNWKRBPpM/deojTqDEOmjgkHysHZDNgUdKcNm8ID907ud9IdQmtU6AUdfh
ZRn2ppomlrnTd1h+YB7GoZDDBjeaFE5+TVen15tdtvLpRnPBwk1eecW8iPST
fi2k8xcH3MqvwITQ0l+hgyAxHKuiTrHq6ErKvAWNuYqxLuoMauEH9Rz/qvAH
dDwahBSSNr6uI5LWx27W+NpU2QeHN1I6UVkweyMq8jdXuZZBnwEttXGJIg0B
2Y+/J8XnQxwvAtstVJgxLkGDzktnHWu7n2Y8DpRMrFNcZUfDIfV8Iqru6Vwe
V9Di48tMq1VanKVwQoqhmZdMMpQcgW4Ew1jyILKCsKitmS8cdmK+jdHa2swX
YHQnECcRCrPwFov1ql3MsToRIisNmOUtGYAdRYZFO42dJGtlXOuYq8RbkTi8
Yo4k5DdbP/spRr5zsYhC9xddquDOf1zmVRkNVbF2Dq6N3CV0cfH+tp4gcFQg
F67WKHXJunvh4PXfdDwwKCfxFHjbOV/HtHHteASufeQPH/lJNxPNNCNxoqVR
jwxcBVXI2apvhKOx/2MkP9yVwG9zCx5101t4rit2+ux5NAp2+F9EQrLtn53X
s6t8D9Ojp4sdRumlO8qXJBljxuJIy4Y18msQQeej4a6tt9w/caNVwoTQYGPj
ypcCab/7OF2XobtB9VtI0FwIUiAVk9wh2RAWghIO8WRerHFJVhIPIaZKcm3A
pLwT+vcyXyKklUijbDKDFjNO5zhjRkPiSZ3nZqNr+vxGAHZBrhjWcyqAXZ10
qluiIuxa0DO6ICc44HJ0k9I2sJUnFtd1ZAA7Txw/hOa1D2f2DNRBtNcyw1ic
QSr5oiBkZEpSK+IXuC5P3kKygldyOUR7/ZXq1EkjX5pOVvyHrDIWN6eRFO+s
4h4yeQKl81b6kO4JJwFzxmaxBTDx9c+4ogMw9QEUfwIwcWaTkvoGXqhB8wjC
KIP8EQIc7hwf8XRkv+DAFaDwEEyyyd02OORT66r55Q4Z0VAOSjeeOo8uQQzU
yJftchpPUTXGZD2juFzbcHaxeP9I07/Pn5E+jP+CBVc7e0+jsvor/LIvoj9e
s5+g703sAWmqIhgIcdpiRKpFtjkqfe2VoIe4CVH7m4GVt92xzwgJWtOpLkrE
vHzc00v6b6HOT7YoVd+fnlFibydOTMWhpwAgJEBA94/ucLg1qgH6LAZI8AGk
Ell9Uzpgu5GeFnHUNJnn9w/jBzYRptlhLAwBWht8bHkUHS+vWcJYf+74X1Lt
0W9z62zFjwrf51SEjvanM3GOqTNGdfjqe6JhlHdUzY+U+UcUQACVFOCyDRSk
50oOvLJRdEjx4cRV6YxhZ0eDksTo5dQUDViZIlGbLwTqlBsZ0iwCDBPIiYlr
LlZgokPm506O6CkwB+/KkAdSG7bh/KSOeM5oDLJ7346LTcM23DJhI4KhcMb6
kSBsOnEJWjAhnX2Dyn6YRTIa8mgsUI7Be+ym26nvffiP+APz+PFnH39LDQvo
U9YiK60aeolVywbbAAaaPzo8O0+rIRffaO5+GSQFJl+f4Dv5Cj4YbHwmQsjR
jwTxKGwlQQpxsP/IDgmMBs/I5JBPSerd4aOKnQ2bzUEpYB+OwBTh6nWT9TKe
D3bE87UUvAgEInaj5FUcyXqMU4H5ly/S/vozZ57gP/GeezL7t8+Q1fjEwcHr
rL5FUachTz9Yp+6P/+RnrzpDhxFz42oySTAI71ktN1BvMSlbk+QIWL6fbV27
hIqYXek0SB4+gMqwTErOmfwtvHmyydfkvoNEfsVbS/0MmpPdVgPZYLeI+0V/
Y8VVDwrJ92kpHOlCORsjkpBla62KCoA5ij8jWkYYPbJyEnaplI3eR9wlhwGY
4i+WGdj1GXkue35fFNCPOD4vuy6MjGiecM5//GsnfMt2+vQVIdVtVakKJ+og
FiQ9tw+q3S7AC3amt19XnIg6/qN62F+ZrKyjp5ratEmzzaV10ROhztuy6V+3
V78BPV9pzFIOSjJFpmrqQYuY9c/ZNAnXE+P5jhVxGowE5QOC2MSugPuKQpET
lwMv38HH4wuLxD83lhNZqSQiYOYBnGw7deWe7kZYp7pPhxO1smgt3+VZStXv
A7r29EGJ/wucBDMXLV9hf2XQmBnsJb6DbWlwrY1+kHmtYvPZOapgKdMrX4iy
xpANeKlpIVDu1VicvV/F6omi+vDoQxbuGysIp9wUwgzW9I3Hgud245Pic1aJ
FwzXqBkpfkXi8t/n930xV++25l9tBD+Q9O8HxwMqDvEDtCLV8hFl7yeQuGS0
BL5mUDT4nW8YpVF7vA4GcyLir9qOwrLL3MS3GlKPkSGhxcROkOMdX08tnjHf
YBoO0lFGnX7r3HbMMy/0CiiY04KHFtGzJu6FiZuSJf9UXaYztPWg3Ce2AjUF
tsnbLvooy3EC8zfkw3UrYdN2bt3sQuHfmgCt/MXCrgj2Epd42/jNmI9LCqtH
/wNgfjinJUQq0Qt/vZkRe55iRFUykM2yhHf6JcBqYflewypcatp0e7hPzjz2
XWZcfvf7GIJ3X6voVtXB3ajQN/tFKjy/H4imbJp0i5RHV8TRSqj+QYJqA4tu
xQ2KW4YxqN3UjQEJPigCcPcVDF3E+EeJ4DO5A5eTJKldnTA/dPKliFYeLn4d
jK+3IN0cEksR6dgGrvJwqd7NxY4kLK3tcdJjuyXT7uIdIDiSJxrkpgm0Kw0B
klY9idOi87e6HdyQPh/1zHimo/3NIt3eiB4vQSUlHa+SVVwjzs4X6bzBkza+
Lehuf9dLWrLVvRqtP+5U5wGG2LKu1y8oJFg6Wkshujr3bZtNp/+iDOBRpsPy
zh00MZjkmIZe4mfUFZ0IKczk90/Tx//5qPYW2muTxN/UFyFm8pJxUit7DudO
AeynpcdEiI+I4L27jtG2I43Y6EgxeuOJH9LP0JQrZiWMyDMrIkoXVKkZve6S
aMs28VGZvlp/L7D6PF3RlopYfKS7d2JGnVI867gHpDsN3jhdH4+gIs+yj2mR
sS/Fy5HrKd+0FO5n33MpEhlnFQVgP5AU8EemN5d0sSUao16JQ6PaaZ6Brvnk
KwtJIIjXxSoW3eAf+YnFZTlUXXwOja9FP5CDAzGyCQMHh/8C1N7rVKNgRle1
FYe1vy67Myv1Z/cETRFzrfmg+NLZsGgGfpKDc+o4svBYHacXifXJR9xR1HZ6
BHYDBHjstViPJPkzUDdslVrNpdrXkK8psKhBwgnox/SyG+RjkEz/xHncxS4M
aLvfZa0Ox00aQJjEA8SkNPUVTyaFFLqvUo2JAm/GGsamCH7O/lqXfxK7iKZw
mxSwXG+IE9nw/ixI5u+g2uH2FlGTjqnjUcNwNZAZJmxTVrLgi63Onr7apnbL
oyh8gQ5N1JsRmz7cFVx33qoHVMZjuuzn48iq0KtneDnOtyO+cqoWwafKZqny
FCHVA6VWtpeiOTOocx9VXacil6+QgX7HNa6OR6Wn9cCmtZfssm3TVVN/T+VZ
n886d5Ki3EwNYia+wcxz8qef+XReGbZth1A4UxMYgLSwLAR1BgONOglbhTke
kpYz6+yfTInQYW0RmruwTvB/Q2wn7Dq/PaQBmXX9P9ue7bd7GqkTILSQujDL
AVPzNQxNmy07ecs8bqaIN7sf57NTmAq/u2PKpX+BkIYrvF+RQga2ZxpKuCs4
gca/fV/9quvSmEGR9aM3Od0sk+qPgPdIBds/GFGwT/Qw6aXI75Ulmm2O+5vL
99eSH9I1D/wu2Aw4/nGpXeOrKX0pCBScn44yNzAlAmFXjN/CtJSxf8Fb+7h2
mAZCHWPAW72srYG+ooX8jqgA5NN22d4INEnJ12VIWWRYfGImEtLr4a7P6Drm
49f4anghUuvEuh4MnbXwh+y8jAmeBxOg3YK+xb+b9OCy5hA1x6bf3I5BaCTK
zeWU6wlNyFdbOz7RMhtG7Bw4Urv8NuVe/OATMjAeBjk3WjvIqYhBf6V1eyqc
V0VahYXFUHTiWWADvJZATwz9ETXtbPztEimI6YtRRuiYM7BIQZPQQgjMWXU9
An0QL/mK4D2PbqQpcGU04+YHR4z3Uf0YK4dCQWeDP9UUjtKV94Po7X4LA3PH
gQ1rWLHwrGumIn3GzJ7oWorJjv0MMOQL21xQbS0YPt0vtbROYLMwOqddNQr7
hgmVgoY/TBsk2cxsH1S4duwBOWw+kpim1yhI3nRzcrrRHf3aFhQ6DJ7EFm8L
ySwWJnURVrIISsOjnmgGkc847uIaeSGBPwE+SCrtlrva0fOAL7cdET+ZR+lY
dLZDeUYdvAVtDnd7b5QYGwWCfUe/ZHlLG88upcvGsFaqXPPxQG/cElqFyROe
mif7R8Z+C8euiR/FeUBuGmKcpqmTXosBK1o846pYkU41xpmLs2TzyZppMtYE
A4KcDQknH/bfgbsFNcLViix0Hd6GJWosHuIrFWrdyT11QBJAlXc3gpCyHika
zdzhY8FNSmc6sR9AZEt53yLVA1YuDXqdfxWfDpY228KjW4pYvFf1tmEcCxWF
Dsy1fzmkSx9kxZIWLkw82ixddFD3hkfKl8j08oEul56PgwZL0lzfngBrSnpG
9Y9pJM7PfCY3xlRwxeKL6x4t4EB+h5jNxlv/ZjGoglWOGtDMdYAp2L4DN7sm
KdPBrYH9YgA4tQfRI0mnE22Er8t3GyejnSPqpnWDwbWJXqgUj7R/iz6Ncixl
T7qFakhm2NAn1qYWRmon/qB/CcjWyiaRdEb8FFjVA7lKPYYZJpkzoB+XJVnl
ipcZ46CYm0xRlmxQcZzWikyMsMQYBNDUkt2ncD+KhapeP36m3JFuWU8jwA3+
1jhPWSNAT81+Z3rKzMOVvHiCBjehqpksN+0KoROemoPCLm31P3LBN97U488L
0TuANWXZfbIcb9XcoFDkT4Mv8UCVGagmA1iSxZzlxdc1MahQgPJpBW6xJSvW
qrKyR3VC485mtb9obh3lP1hq/o+5/R6hIWVJzzRGv1DJFOQBaK2sr7+pU/0d
HD5onoP3Azc1NvHQqSY/ArUXkTXlUxLA6WeY0GymwRafrWlUIze71iAKBQh5
6EPfnTOb6pXYjsOc7cBFKAvj8CMRSuwWw5KxMRsdlNmRLLKHARU6lDHfRUzh
ghMSvxpnDSKa11BcR9ffHmcvrvr32quCaVjqNyIfm1YuwbgxV15O1dEmQtKg
eHgJpaC4hTuuPZzNq0gExs1RwcAPBH8MlIJA2wiq7nWn6ZufHfzQztw1P1pl
UezIN1WXvP4yveEi2qh9y5YeJ590xjeyrKuYZ1T7C/AktbZU0nUngWrKn0s6
S1B/Bb6KDjyFJXhO2APEzbwYY1QhtjXeQjaWn5vqyUdkLGupAO78/hUHVZpc
aHa+ciuh2OvQb/SvioEKkwtAgg3+M7w3Jh4uC7zX4QTz6e6JrwtndNpwQkT9
VPsk21PnE+YS7n+Xce4eDwgDT0VgGJdscCQFjjUgGJxOtocDehlXUvQY0pP0
VxOlakZ8450qBQNm6+pyFcFcsFUtlbG6AHaxF+wWvkGPngwRBVUCzi1ZrkUl
LXZzXYvWlD6pv3Kgf8lf8Swor7Jre/K8eLhgr5OnZeUh0ggc/Rhc6Hud9uGF
/jc8NJSuG1EPmu4CVNknoNIZeZlz4OMsTsudU/OqfAYKF2NJCFo30GEDDY3l
AVb3C7Sl8FhrGCsgiJHj/ZJduDPHSsROxoox4Xyi7CcodkuDb3A629yXhmWW
K2evSB8pgXKFFS3IYTDZxd/81xWbNJst+rl7MQqv0PC21H5Xx+VAsv9Io803
+fHMmAcA7TtMKXP8e8g8/o8p4F+VGs1bZ+QnfbIAkvm0GdfmyzD4F6cqlNqN
EFjt8iAJPTZ/aq9HizRts6wahgR9tCfR1LtGBzXB0T43AO+b2wUOfymGACRn
6RkWa+ljt868syg/BNYEpnhCtOv2GdiAkAzk6wjw+VLJ2+S/EsuBw2ACmzze
cQ61jdbkxUpBVfPhURVR9dnlP1q/w5/J6XOfWCmGE4IzMLFi1UBlD1LwPx1n
3m0XciBs/yGNfqlVPtHtywORpONpUsulnqu2GMB7MTJSyVrCrbA2TFWCcZbA
4rRc4j1wBs8tbS8OrpxLlTfHwhxi2Smkrm6h9FHfEMQ2m2HZTk2vEa21mvp0
AhDNnNS3meAhMU38DnBFRt8juqZTt6vz13DsWT4YLaVWjlVTACkabxVbpCHi
mopSlUGnhvugA8rc7OadjPFLRM1DRFKdIHPDGUv76S6gDWXRAEvA4YCaOpbr
hmX6XvEuFW9H90cHjaOG2PBIWt98mDhed/R4H7TfvlOnkUTJQzz/SECEcX9E
VQSJOjTjxVscTZfMIOPFOSVPpSv1VeEEwWTwDVNrg9orI+3FdIeV3Hn00Gpo
7SMnEa2VmKfzuaJkq0CUixCpmdKEFvpjzqWvVSWtqvL0dKwWljnQLHt6pySy
+AECHCSqytSK59XtLW+AyYsJ92F2yT/9uEyVfXp1hZTNTnBQckLTX81E7Osk
V66Roxr8z0uCZfTG1UYo8qJs6C3emfv9EHFqKGV1iThi/d32yPdUyh76xLMi
xt5szzrBcG7bvxY/HeHwO4gti9NnmSbwMXCFDcphZnSlS+PZ9dupC4D8pFHW
FKWUD+OrU4td1XfrBAUcuGziE0ill46gEEJqeUsPvn6QMY1P9h+diuGezGFC
uZsLlW3PoJTG7zzykE8qrabotbeJZchi9AEMQdkjXtIA6tw3KJsowbe6pxGt
YROFArmb/BfmxvPPZvCGaN8yfWwjXn5RT2wA/ReyzAALGl3hylsQjUDfMm6v
1INXRQakdQ9Kxcsox8URKZJZFqUeCdowmkZ5sSAnpPGCxt4lqQmHYww2JnhL
BpImdnLYQs3q2WHg+HaShd0rV2aH4sR+PzHeB0W6yUKjYtdfdkmB/JTQTOyP
gnOBpzncnhX4jNgKcAy2zrVi/yX2gFjedbJQ8G2pwhnL72Cm6dtEejTeyIJE
MA2/Mi0gk09OvZXA3x5O86R7YiKbMzDrpr+DVnkYAs4XauXD3IHrYhEb34j4
SK+5GlIQtuaRp5tyWKhlfWfjm5oksRmiDKZMND2d6LFSAvqKTFeTaIrGIysj
5KvZWcgmbXW0ddMP2b6E+CQzseXKlM/sto1Q3v90lmRwgQ8t9NyASe4pFs7c
dzjYXN4p2CnHgMAjJrADRHrJ817+d+xR5UvvsibTsnVP0rEpc6pZcyE5FOxs
LIb0/i4At1bLdwQMBdMra/UMQEq+B3XpUxWgQ0XgLrRPrRfcIAwQoeGwRfpU
NUmggymNE+0b8MjGxYDluRx6FeNJhtqCCHyhN9kz2ZCwydIOFLgaCke5eRW6
labaZZacWOolgxp6tAOEWov6gMCsKAllHWfL3AMM7woe3Xm1bBwBkWyeDN6U
Spt7VR2DfPN55g9EFD1BT9xGxeuMCjfmffu7coMIlqiYq9Svfy9OFr3qS2bM
WbGerCVSSR3BxgW+E3pJ7FRzhL1LzAjuwJXYx1XneBvjqSH3mLLhm2VSXvOV
ARb4rsubaVBI9+OyAn/FZAP6Or7mAiw3U44YLBlzBRT6H6YZkwBlJvYCjveG
mXallHezH1WEnolZHnHMJmoTbu3Z6u7sQyounATEpLc8uzn0l/WCSNtV6ViK
k89/FdZZUEpeWX+xo0PwYSr05PfajmLXapT7Ln8dRYcqGsFuSya5qYr/v7dm
uv5OuMfL5g6Ln0eL/1FKgz0vPBQKCq7BFYPyAUYe5tYKq4dnYwKK5TP9NKHX
VqMipBpq3F3kTIn8/v+YbWBgVI8MmSGhQDDQEyszsQiMCsQiu/5ZcSBoI7qN
qOBss3O4r+9ZgTZNtglp9qSx9Ewv773tM2ciEjreFahAl84VAJsCCh0It/0t
3BW1LGRDO+kEW5JgBTdwnagXbkd0ZOVvKCQw1/d0aIhDawq2jezTfUAuiyhM
Mljx6jASOSZK3eodbL3J5Ly1SFrSSfXx52Uu9zKaR2MoIZ0rQSAPvwwasoe2
hphrUanSswWlH38sW+7wjxsB8zP7amvWbgli+xczpZo9Ubb3txVgwEICearg
2jgTWEbqxh7bR2p3e6uyb1N9AbVVU3mWkD9sgkHbtwHdNJ2IhmcSxSwrprnJ
hdxQCY9MfjGIpvpJiRYLaO9z4x+1/htstg9P1agXq3M86dd5ZvxQcxodMi+a
bq4L1iUqLXs+88WyZgUWXbEeJta9xzwl5wkiQ5+o1h0ElL3921+Xuo5Q0Mbq
aB16/MO6W+N8UvzsedYX5ThuoG1/lf2tRPr7rBFjY8huVHgrmNuy05ZBFkfW
60I/kRvi8nXn2x/wmMK7Q5/M2GvjYW1lkhRxoX3x1dwxxeiqbgX9q5MsatUF
0GtgJ388JAWdjixVZYPoI3SLkQHMx0HGCiLMlqH8c3G3h9MQVrkhvBxbeqFg
qRn068LX9mjS5nr/061UmWISWtiZqlzgKieECVheqvfEyG+soEzv99xjMmUm
MBzR28i2sOglSSGRkb8KajO+hw1YjyrwURZqKPIukJRy2KcaD7Ww/dQ1MT4R
Pf/ci72OJdIU6NZq+A1M31LP1TuXQfL1BCxgB1DkWZNm7lWfcr2/aFICqm7Z
QKAIl9fk0ZEBml05QH9nVovB8wdq60Z4Ay1uzzjGSfRkVPhS199m46Ax/0H2
gyqXYLlSBf5ThvulpCBeWSGq1hJC9faRU/XHMusTL84ufBZsan3+83/rHrI1
gh/ynj6EucDN85Vuw6LHoXTpuMRd7P1Hx7kacWEXcigIuJfJiBHSEucpKZTs
sxCE5MjBwum5lkqJTAfoY+uLU8uBlG1ZQGjIvInt/J3Lo0ySog3PCd6YIw2g
2XEUYydjy7VQrrsR23d3Lcc0tbwdAX78ZXlHSHaDIZSgyiiDEC0B40rz4iTn
I/ESTxtYgg4Dzlw3IsG5PVjVdCYTIgN3Xxdze9m3vpsT2jCybdqXrj6PRHjW
5JRSzdz1lhsUHiPuvyJ3UY5Xgf0p6M9EuceFhZNgakg6JVTVP8OMzbOSI5Uf
V+ewvcJleDEvq3OS0NJ4c6dq7SrN6BnXwZZIY3Syx1hJHq8v7WGef85wIctw
E1bHqDb74wKQ9lPwoEObhzEIY0UoLCJcff9IWjHwE9Wjqbk/DOYkfBVe8yCQ
p8njM1bgoijcz1Lp+01OFMNw4iBjLWhY9XjKFqKtLDq9mwS81quh+fKcTPtE
8uC7lzmzUxagpLgqbpjM4RA2UfNqlNReAWOvYGqjwn+deRLByg04Io4DBJFX
coZqyU7W5hHd/doYJTUzQlV/7kIJpc5eeLB0mMOF/W8uCkCs3vISDlgwyizA
eNOSWWnRUuhFqzEcev5ZLxLHGymyY9FJGyujrk0SitFD+moo/0vpojiXT6hP
4aD7wMiL9cA4kX8MAZBHy3oljFq5hjyTtEkbbkpWdt49DRePx/h6fWb7PlO/
sPpEHXEwGC4mrBdIFm+t1c1XnxdAXfj9jQyW2XLGPx4x1rsNeFhE0Z9jsxYc
tUEwHdCxEVh7aGVN5I4t9bMifiO8MGMStq1cr/1Xqyby4jIB9j/letVnSgV2
tyfaEkofRhgq0o3isw+AYj2oT+D6vgrRzIX+G4P2oz8sQ+bcdLmLjoptGXwi
FeLRe27Y6j746DA6ERo9hLAgYTmmsm4/F1BLyN2fKwvBYCKIH2aprpQDT0B8
NpyJ47KO9GaWnLoNL8ynnN8PMhLZojdePOLsaEEokJnUMCiC3FkRbK5vddYa
66/5PB6ECU9Y0y0RukhmLO/5VVQrC9KoP9jhDVKQtF5XYb/o6k/169A3fOqt
K4zp2OQAjG7jazGJELT67rsQ1EGoi7GAfefS3bo2jFxpfY0meXOhpvjJGBzy
oqv8MMVg1cLoojIz83V2JxgyvblPFUTh5Haf7UTeR//h/mEib9UNPv0ldIvg
tg4vxrkYjAwEO2aKjae9dj3cY39YLfkT008no16q0ZrUn9iq4ypX8arA83JD
01dMEZ56JTplf5bO9iwHj/21NoxL7zeYkXR8Hn9vqqb7kI3Evg/YZB7TIM+s
JyNKIrlkWq2rwUQxgQHYNfWwC6LNJDPTAEQ2lI0kcFdztJXolLO7L6DwGI/i
d6mRva2nAGCKP0tZg1OLHLSnstB2raFHn/SVjAj1KWj+vRsbIVyfP1aWbo5e
jDnEoVFFzZ2BMphsKhNNXV4oXBUNwk39kDRr9JYerCrE4jc7ikw3TwmH8jNE
kXcpySNrczfOLcG5keiyVURqehcrlUXQzpIrLSJg9WObdKr/YEmmm8A5uKjs
i4VSMQqnoPV/gaGUwjxhTuYztdfMIQA+2G728C9A8yjCDIIy5YYooEwcSbuV
pdjbUs6PDI1ly4JRYz1b4Yx73v3yONFwQ5y8LgLPZhxQpZuN87B5jcnqaL+3
PbO86MtfAPkrXs+T+auma8x7V7vqz1x/mnZ9LaTaoCY9QQuGRqjujuY97oP0
AsWrJwgGreCtrQzcjgH/DfHLD3EFKDP9KScqdU0uUhi9MHC0BoCrRot4hz19
g6MbOr73AUnDzXmq7te+NU0A4VwFYCrgrdDMJGs9uwtJq6gIVyt+cUxuYihx
EOmX+BoE/4r5lIaLH9U3wihyI7OsPtKnGc9IRuAl/k2B2xuOlg5aC8ahMwea
AiH5hq3zjFvNzEVuwZ8+8gwmkiQrL6k7J+w+eZ+QvAeBntAhnZmJpjV/y3GP
V5JyF1U1gFMllDBNRTsmlwhxHrrr0wI7L3bq1XVA2ecR6F4iRDVSGWJgHH82
IiGJGFCptNAzbHUXQWj/Nd4i6as+P4ItiwSbRUIsJjEyirMxqELfKzag9UUF
4/UD4r1t7nyeaj9vp7t+/Q8IRaREeujhGZe+7H13U/0qecJQ0qOYoDVdWZlT
wc/lpgUbX2f8ftLxsOPmaz7u3ntbM4ZoWdOExvWmvqmjqDYt3z5zNy0WwhCd
wWURu8P1dMd405yTk1OcbqEWEMPtZMmQgU8Zl8F0/cGWMIuIqhCF1rQWylNy
VkumKlMoKkJymJxBGVpGYSB0d5Afxuq2xqxSMc7b9aJMp0J3KnTZeFEcqVjY
Tba7X1ZztnkFkDpwpqEddAAvK6CqOW3CL0r4pZFxETCBDyknPgqPJq5KM9y8
09R3/zgw4i0PAGm4k+XuzOsXaYWQqU3brRfoEK9Ptu7o6PsKiAZa+hLtJHjg
1Rd34DBpQ01jXNPVymHKzfmX9kFlRda5Scl+fyMHTBPhNNvSHBzQ1cHo1Onn
xpClHcvgqAWrKJ5CkI2v6j06RKJn0Hud5oOdO89a0uhio2rq158KYDtB6F5M
kYYmpYhNtG1LK+DL9yUhhzy2I0M/nGjgPbnkxmVFsQjATz7zL8nAsouUD5nA
T5MqhgNpp0PaA34XGeic5Mp6ygY5X8XKL0Azb9PFnHkNQlaWyNyGAwKkZSKb
JlYr7ANrTYDEqGhmoYs+cQ0WP9nZMNu+3bbeFPkMmpFa65I2HDt9QBdp5nn7
Shu5aN8diCAtCP6+3zGC8YvJezGQ+Y6zDcszeiOL0faZKZ/WaFfRCVTeGWxT
niWHxINomWCTWHGivZxRq72N6wRSRb4xmlPTAoDQ5/wP9tToV2vu1neaJskM
tv/A1xEGO1aKbpWGnYVqox+Vlaegna5RyLz2sdtqlmgIto0bBlCBsix20a2B
W4Ojez6wUqiQyIXvN7c7VXA9vfqrnFtrCV7E1x9l12txYiSrk1OAusLrxuzl
T5priu6gQX77gRF9aavguVpY5IoBN+ZwTNPVhaIGi0aJrq9ODa8AI/8D1NQ8
aputUFTQoWqcoXW3q3n3nhJpfxjXqt/CesnxKf7qTr2QnjhwKLUlob5U+YPp
DSa+4w6fFWHsyaGKw4OZNhoDWluZXwl2WBzyfJOkDpIbs9IYecNQaHc/CIYK
HT4GcuQkOa61Mj7y2mGz3q+KrKdCtuv0H/IWzws/kfx52N5yS9jgEZQ3/t9Z
SqmqGTb4tlHpsR9S2PnnysJds5TiunFQ8QVeKrdLoccUla2hw/afJeRaJehG
b5MY7+VBtFM2qhcIuD0vwPrsdHT2AEpY1lnsWBpsF8Uq5OIWKQxWWSsf512n
MBYnUOXEsD+zKZGPEGxaAUjOexi3ciLrN1Acp9TIi1aRw39Yxbu+JVMFXX/Z
pzMDJrEhlcsChKTcEdY4ZIJVzeRPvxB/iDOgAxYAu2H3twHk7SP8l/zIMces
Y0qki8Xi101270dD1ZJTxKdh1PEemlUjaKA0BdC2HTpeMv3gggzqd8nm/5/1
PVWGOfBOeMa5vV/UGt+GMNeMDL5f2bnfRiFaAVaQbZHRnNMR+kLCMMv3mgJZ
emzHGQ44Jfi8E1m7RcplbXKpBhSVAwP6zlbOM/3Nvkbr/h9J7QM6fIYapaRb
kXKEHvKDnLDnwWXXkNFAYEbRkrX/0jh+ZER+FHRcngIKA+60NKN4E9rg9EaZ
rPiOLsuOI/0Nhid3hRTUDgpyLk+gahZJECK6oI/cRS8FPxnn8TNHKZhWwtKa
tocjslvxqB6/48ginOyW0AzIlzqWuX5haa+uMJvvYlwJBA3BF9kB+d7X9tci
aITHZ1P2+xd12OU6gnGEeOM05ElcFjySotKM3JPIL2HPIA6TasI9Rt9XPz/3
VjQn0xGAUdq4lW6DZTHW+Dikj0Nn6Nnr+R0GV2PNAcVSnwQ2XQkVY9Wh38qu
Flw/Qn8wwj3zmsDqijt8wMWVYuwqhR5atP5WsXxnsDVKJFz6PhElgQj9tGMD
bSUP2lesIfChCKFJ//VaARbuX0af3qh8sb7+6Rz6j5KeBK3QYS8FlXOV5N9e
Vk3KX8ZvDDmUK2txgfsl8ayl4SkxOXvfemjYllFbh0nLP1Nx6JcKfchaX2bg
UlRXS32YJ171MI59yhHBz/wxj/h1O2ljWRUHxSbMUpK2voe3s0lSyrz/jYJI
xV96tI7tEf448492i84dm0ovB3YwN33tjs+CAmX5A4SAsm6EX6jMfrg2e3/x
MY5d/9mgZeW2zvTx7+KrPoAemBC6P0tShp6FJDRkpDkxxf24rhiO2fH3LX9H
xtVCrPK7yQ7XSq+YSA7X5gnBvSLPTvvTvaR0SzYPTZgK7u5dXxh8kiY5x4DS
5U3sLRZgc6vpmJQRcvQFVuOkti9REUb06NENTaxoLaJ7T4AwXD50MXE0EdVL
kfkZ0pt/RYyWqIbJVn9S9aVo66sP4ZnPywp6uvTRvBE7My/T+2tbtMiF6JAG
WQjt9EjiDTWWoyxZWoA2HzbgooCX3HCzj8bBr+7VoKKpCmJtYJVRLHZwiGT0
Oi4ZchqPBvGAQh4N024U2PjxTV8R7F6JD8MRk+CTzklXbLLcE+p5X3IQfOK8
9U/Xnhs+f9H3locfjtQP/kT+VVDCM6ZHW9YQPAh+17a9jetp+tuRU08jPFu8
RHdXSOofoZfWjxSu8lz+C6qDEAHsIUUV0G/GtUOkRFZ4K9s5PwYK8zWuTUgS
oQFwJ0wkJGKLfp+DNzM2sx6Mu8YiZr6F+/8KPbze5C4656vPNoTaVX+kriOk
hbIuDQoOHNeUHWRJIDKgoAZBENzdeaAVCdShyNCI4F44RczXVKxNtBENDD0z
E4OZoQPvFeyAscOC1hXIzq6i6rEFms6VfAvbBiIh4ZXr0A7Q9hVdu8I6+K2F
SeYBhYBkTlvLXIRFnLhIUuw0H1xUamwQF6fDaBEFD0sRUs2YxJ4wi9Jv6K4p
5ILgxwXICrlc4PWFsoXuuSjDzRxjYhacxVjKqbZ6VdYuahYvZdsfRnZBgQNw
MMNvC7Uu4BNBlJ2xF+E9lrGMuKL2BWKCNxRaw2RAmxc4e0wz8Xuvx05vT3RY
Vrcy+E3JvKHBb9XbowF3lLPDC9B4bfhjCnjSnL5J0h9pTFuo+LT2lTSpDv8X
vGQ0Xfj9vCEg7kj/CqHwlBnJk+YwT64rIaVn3gY6uN0Op9ggDHphLrDmvU9x
HWGdOEOm8C2KgaYwwUszUtKtYbQzj6tAtKIY+xFgYotw/bLhs4wXsVueyrlH
g2LKDAkM0b7BDtXfqL4Ef5L4tO8lTD0/eRbQ8dFJuLh5LAM4u9EIss9B9xNG
wfYgU3PEA0wDKaA6JhSHBPUO+fWOX6cuJcCsHS7hFEYkG0JTCLUuBxgUlUir
GAkYJFKipkOc0puiBB61UzDBISZYLrSaS36XBojwwELBcb0FvMF4XcMSdwX3
KU5WnB2C4i15FKi8YNp1UWY/kxsihFkrsvKJEg5XBzSbAHSlXgBrDygY4U68
Vnb8VeKc2Z+vOVDdVghR3dbp6auAjz8q1USrPjdpuCWmWoXFJU4SOlyefNZT
TM97MjiZTnXPEEDMkJtbmSXvyE7DJQHjQy3Yxma9x4pnsD1zAFSxOYP+nNVQ
9Fe5NFqW/YO+bGnu+93kqLqzj0jbLPRmsuj0QUCwU4IUx+Yj36ERlhh1NV4z
KoizDqLbA21/5ADJ8YZ5Dthm3br/PMP5ooCGoCI4gkzd6Kkg6jtHSi0LuxB3
p06nGIecpWFpnVVgcgGhpvHJ55mbITt9lhJFVJvn2AYydggz8AnwQqkstI/b
kwrZ1PRxKnPaqVsrDl3Vs/BNR47oxDgBDkmQwMx/a6Jr7Ep92PdpwR041khp
V+tmTjLP7KGEw3vWaFdSmdf+0YlmAtMCa7qzyE4917JBggoNk7QIpLM2mlVc
e4T8gBImq3fJplccSCJCezf0tqWmBkk9DSBWE8GgC8zmMDcVR7KDIJfbNhaB
gFbnLP3Qt46RsB+qKXtdz4y7fq+UMajZ9Up6xXbpU3TxYrmtt/81tshI2Tri
y+hVYb8Sa9bU1jh9oWAmR829/P/kSAbMQaMHLZd3ndn/7fYU1t7SLbte9J/4
ageE6aINDGT1mW9C2Zl+Qt/3OY77D91OhZFXOwtoaJfEnLUzxZTZCHRPLi5J
sXBHSWk8ux6T8WsAdx5R/w3hOjGE6eAYi5RryW+yAhNTHYDURvF161MblWrf
DnZRfH2wPBc0bvam5Hdkq8DPHElAeY1hEsKoaHgHJ0tJyenWSELqSfFIbX5K
RfQOezujGvX1O/iaMpPB49TRGpTDz6OoICIeMuvO14aWNeLa2k2D+CY5lIeb
Hx4bGmyyFQyRbxpYRYJDwyaUf5YW259CB210sr5lmkyFb1Vi6dLY47eEh0Wk
/Xs40SeMEm4qqpBb119cZItc11WVtgryTY+pEoXZJ3OtDobetQswiMkPjycA
kH7hRyCYM/4wGrCDLSkeSVb2SP5BfpVMHaLV9uIEOSkBwNovFs1nzx6b2KEe
n+zjjuo65WeqZWYzP2VGqF4KK6jf7xIE6ggy859FCcPeMRcazoRNTehJXU75
n6rIWspaBsfWEktb8TqCXIxekkYVYLbcdzdPv7EAlCqaiSKGbDZO398VxeWI
WcFL+0vm62zFRNkdD9FhDjvm6rKWM9qPb9t1fQ81KdjQA4v9r3wZ/ZKsw3Cy
GWByvV/Y0bwBSKZVapiufQu0ldylsO8IAGjdAfeb6bCM9VW/7+v2ORKQ1/Tb
J+8of7xeXY4dohZ4pgXaVbaPXIdanPtp6byqSUB+15YhIvMryUn8KnI780Wd
h+oAAAO4BQr92bNkeTH5zGIQ9o6zEVz5W50XIQW15K3fD4XuODILw6tEOSdC
HBIwBbg6EPDrM+mm75cGaRMSBZ/mceLhX4wL2uvmspuK8KppSiNfrgNIDjsQ
PQqDJax97MKOFe6WXfNfSunOpDneyD5VpO1cpZ872cCP2O9Ejsbwk8Eaj4Xs
WYvgcRW9wHuMbHkI9gapigKErGjVHtLOvz+7pwRjD3qr+a3K9IJaxl3+lT5P
DpII5Suqf8dUKNKsOtH4chMEYJpglpLCfBbxdArQI42ZG0s3khVk8lXq8jlZ
7a/pGKwKSQTRpuE5YLkAr05zdTxhJ1gT139w0qozpD0ZsAIep4u/PlMhYFDO
GMfZT/lH0EUeW3l+EFPpY/ShAMfoY/ukHih2jhJpsOuzEoQaRt/99gOCf025
8uMOgPcfjJ6oUOmbrx7RgNE5NVjALkFhfWvxicPf7d5pfFlrkcCzu/hrh48A
vz6esxbVhIkvBjeaONyeAgOnhvvKOFkInV83I1NgM2mzQr9/vJgCGpZuNvga
CPb8Dp5u3WAomkfHzIjibjITUKgDPa8qXFaru6skRYNhGLLZIFQbtDDG17IH
bfYLVIiKni/jF+Ok0CsmqM+X+TMWp+x+AkTJnBY3htBY85CrQkcz29+0QyQo
wyaW2LcRNwHuBUWRHiaUYUQOG7PacUlyuC/AdxLWo9+QnP3kPWGZuYubD5En
LIFkxyGE0lfzde77xuFthCSoidkrL2B3e0MP/mBiLBaxTTM/FdW9ZZWBhhER
I575ScZkh9ruOwwFR02TTGPZcYVPP9/vIJ9bMbuNHcfDJoWcEbIqU71s9Zga
tmTXn8QqiM+lWKUcU/Lm0g/uqLhpnfNEVPBSXUDtDw1CqFErhWl1916jrqu2
8o0Xr1sc+HjPq96KTwO6EyKYJW4Ki7rOiFUPOXUjxbHLTm0T3O8AOTzBqzNE
QBgCUhgj1EcIO+oOJEnYa41jJq8nlxNaXAwKlx799H+RoK4dmQ+vxhx+WOoU
eP2d7W8ZnMsyyWuHGxkmh8uA3qnm6ta/edra2XVKKYa7Mt1biuq++njdW/We
GJouADS+IbLMzTLnUmkWQ0kjTnqXwBc+gw+xzztaQGrF4z2RWLcy029VZpgY
9Y/q3txTyiNpSMg6gDtI1zqKDCWYnlucSOxsdltjNEnkYl2aQ2S6LxANGYnq
/JEAIE/a6Pyh3fnYk0j49JthHJH+531Kgk3ZPEQv0j76moYWxpmCAxbuPGrB
hPqUty7zWLU1GcU2zaS4AuIVggR3pHlCEE1dBmyxsexveTDsTuYT10PGNGrG
mPux+bo321o8KOO7lIh+FmACT84/xWBOsSs256kA0reXehxHcawDerpDh4im
a701YDfy/QtBv3ySMS67DRgpyZ8IknHB3lWykPvzb1qYcXVy7hTy5OxjJm++
osCy1nN8P2wkVgXT5LLv7wpUR9EPVpNGQyv3t/iZiIf05YTm0EcCAUIv4qFI
ui56eBGAtbcrZJkGhFinyw31EOf1pN/k5K4OZeCUaIM/W+okaGjHpaE+V7Jy
qt7doVZs2h9CAcCFaT4WBYsVrgpWF7T/mLMCQRJdV7NXzZQ4SO/t+3d5metC
r/qcr4w+h0uProKVthPTPo6mG75ffUu9Fnt7c9310BMfu57cWTWHsHT2rPHT
wEBhjWDki3pWKz+0BkdVFm2iMVNsoBCeWO2eQfwxsKPp67X+r1ToZMYzdNNE
MGTZWKpYLk6pr4Bfo7wMgD8zPAMGl7LuWyl3VncXQzJknNdgZ+nKeWfnPfnU
O2E9qJ+OJIkjIToZrOcTxJiL3PSrJie4I/W5U/TB8WVhMlDmJvVIUP8iDNLy
2S0IA8GD61y6NBD0FXDEybQ7bYkzRsATSHVavE2P73ITqgwT9e8/EzOOmmtS
8rzUklaHwyUS1IIGQn5Xy3wPmLNRnmzTTLO+tujveaVK4aYamt6R5cGUZwty
7mXkKuufBkZsbxU8+RmNPQX6KmcKKVHF1IGfVjhQQKejHxqZ5EpG38f6VKCc
gB6DwtPSwv7R0b8aVwpeSj5O0tdavyCqmKcD+1iwV6OytsY82r78GZjk13K6
cu6/rlK+HJ2TMdc52FTSJ7sjBMQ39M9G809LAOFEfrkS+ChNcaUcnjA3s8ED
seUoj5IblStrg0yPCxYR45ePm+XhWKYCfvlVZJ8Qjvzzv7EVap1RL4jyzdu5
w40+pmTlP5UGhmy+/vN2SnqcegqtEC1CwLbTIsjn1rFan7dmAvxGKjSNGwWK
9m8nqJ+B0c7pirGRIbH/GtCxr2wQ0k3hmzRayWCaccuVlU1LoclGaLd9nVZH
sYSUeC83TvzWS6t3u1Oo7+G90AFQvwez2L88lc1RX0h8gOsvaecKSU1AurKJ
tK1JF84Ru6CBFJTL/5kwU6nGGXIwzmu6y00H66/J18aRd61QoTCWHNbigk7X
ViDcMJw/iyjqFCqm4ja1L2WxAhD0Ldoe/5bSvqg91eL6u3+Vrtyg6486l4DP
p/EYvD39WYG07ZoZ3wpcQTobu9xZDSD8VWvEcbFjMNYL81FlKpiMHmQPvJGL
73Gf/AqxTj/F/GGha3UrWqaY7a+b2GPAVGgEb5zpo43lykm7qEzYZ7B1iu+X
SeCUKxIy9lESNGj4SwpRM+HsB1HkFhz/vCS7kTu8N2Ye/Afdm/ynnBki8en2
wh0iksnbs3wFAbdK/f61KUBYxfWr+DANvCNtY62DveU8qxsPH5O3q2kuqJbX
0TrKVt7oUaCdILci1mKGAYryHATnjfe2lb15ddssIGQHc0H+7gSp/w8GQ6AH
IStlXxmNyj60MnSxyG4Ul/9l2Mv3WgNxYlV29QzQQv3gwbf0EOFfJU2GjEfs
vosbBYAzU3LS9J5VpvAkci+jOq63u2CBNky4cYbakx/jsBnOABrhRojRXzmC
tNjwCy3xRHSsAoABMn8W58t880YQkdqcvMq36rjmYBJmZepsHGRcUsf8xB9h
/h5XuI+7g3Sh14qYE0EWyzYHZ/hhr9sSito9wGKT6ih5fqZa3Zt8sU18hhLl
1qUIOMgnzd9iC6LZq4T6WBxWc1p9zU3ger87SJI4zpQ13QdGi1tZvJajFqVB
VqvhwNHE4d3cIWh0xrGLUOqgfOz0zWYCjnwDmjKZaM7CmXVSggTcWHaQAtwk
mtwswMLSY3bYYU3a+e28u5jBx6ZhDrS22zQEkMOIj9Qd3CV0nEiDqkoGjerp
6RwDBXu4y8Z9ogAlIv/PQkQuax37zbSihioS6k6BbiJKV+1fz+zVpeIrYX9s
lDZ8NYOj2aeB6huRkV++fXvCD+tP5Hfq/tZBxyQalWlR8ojV5eLxdB5dzE2L
DH6JH033RM0NmpJ2z6avRtuQofX53dikKEvXLJYnWylGU4Y22FWUR0eSH8t/
2zsxDlWOXoj+hS6g8bEDSzg3cSWbu4MtQXWStn5d5ZN0QmbTusHrAJ1NQr9/
F3F+rsBo/jnD3sWm82j/KGEmQZFF1OC/efm1c5b1z6XE/uggnCPELp/L6od9
IZiBSXsBwbiU1r4dLBhKm8AYz0zV84R2kBC9gOpNJmRnOZBwomZHelvFBEbE
zgFilElYHQrV+3g2Z/03o0UjkQe69prFviJ7dp1PowFIlrdblDw4/0BRvQ+Z
UYaA4VTFIlxr72nUFNHw2qRhU+UeT4eLBH0aDgeagxJGlFu4zkS/333usgqZ
PWUO1cZMFLUD8cBxpqXHYZdFWxk2k0WhzNwLpG6lsZxlf9aFZaPQZQIqw5iI
mz4xAP4FelVD3/JnMeNz6lzpoFSx7xhgxgnZASodQmPOTw6X6vT136z5mbKl
PsQ2UwkBo/2GIp0VRmu8q+kocJoQ06/lUGZlWgsLFIz9MPduuromR+2ZRvx8
nFu4sI+wYmlA8RexRdqGj5XT946alQQlU2cA+usNCfASu8pt6qrdtL/HskkH
o9nheNwWNAltTD62ScKK25f5sauvTK2yz22ek3ZO0msixcA70rZ4UnnNG9vs
pj/vr/8zjfgwXop0lG+FXTBYT2Q+GZgYCNgJXMkG2qsjLhJugvi/oxGVEbnj
0/9AkzccaxdNlLIL4VsN12ha5sZleAmdsGuuZBCfAGnoxYeuiPsl+IFrO3AG
7K39A7kOVJHCDuAMS8KB5S8BNA5qCArRZJ23BgBpYYuO5wMi2l3UExGTmXpA
0Xzp24BuHQv6E2+CgC9OUQYVgyGAXU8TfQoX5qCRYhZKnnhSVI4P1d/RMZA1
D03Xw5c3aLg+DgssZRMCG6/i4XbOM1pABzV0GsRTZERSRQ3dqtJeOw92fxfj
Nmize/I21WLZwS1DrmDTQWWGZG+BUHUiKnswtuz5KJV2X5vVlJ9jGZI5c6B8
wMIfu2soYPcyqDuStojQFTuI1lXWkwVa10KDRD/svdKUlQw7WCvsw1WzQp5R
wnsqy16odeacHIYSFg1cFEgxMSObfJQcUU/qOAClgxKGjzXL8kXAC2HUFhj6
iyjtDLkLeVILt0mF++MaeofmiimFgYnciRS/f9mi1Cj8wVCNBg0f3OJSJrUe
QOb0BPmZH/BGoeL0iYLdNewbp1BlfDab6lDHjClKl/YaIdyEGouFewnO3JxU
E03Oz9k5DXt/Y1weCZJWBjQkmOauFwtUFYfcdgyNAPtiO9ri55Y8p6O+yPz5
wG5UO7aXklDbMA9YKPvxfxzfpjQJ86sWhe9R6h4g4Q44b8vg5NUBxmpGpY3g
5x9aoUU6zkzxT9HhR1IZaeL8e5Embh7ad7JD77SFcLBOOWdzbmfmburBTEja
gI4uo9N7beXkAytXIcA+Jl5CPzmZdAwUfPOxRHhk0eKj3FADUQNEOBE1BBnK
5kjf8soH/gpf+Dc/nz3ZuP3AxBzoM7hfjAumCwtZho7URwn5eBoAocR8Wy6I
RuRFiiV3d0jkxXA1eahq0fAOkWwJhkhPwC6SH9A//r+WRK3IAIBKx13X0A/E
KK4M0iiLU97FC50wAOhVPPeHvef0LQRApf2OjgVS9tcHMZMzIDgHWGjrLHOL
bi9xDE5X1ibFTw71mTPUHUabo1VrfYfvm9Vkr48y1t/7Svrrh8VLru/UxV3x
22lqeDr2ovw4WTEkb/nAF1LJfvkRNZb+ywwTybRzxJN2MrRpJgOskc8mndHW
l6XL2wOMyYU2sLHeLDW/GBon0f+nkT0GIjY9pQxZNTU/7tpR4psHUsJ0hO5q
nDmQ88BRIOId69TObYyyi7xJy5wkdvf3oHWqON7srOEPJuJYoZPato3XuHT6
IqIRKcuOg3+RICHwqI/+5ddSLgs6tXIgKg5OVh/A10hgXHuSwkAxtdp3//ie
IL+4RrffLOUb614TEClizeOWXz7IZOkxqGcNeOjh+Xn42MekGa1A+lU1u7Gu
vpD8Nfrs8jyU2z6WwyO54WX6jkK5p9QqwNeUdG4XQz4hDs9ya4W4ZgdwGJBh
IUpInOW0UiaOlOBDoFQzD4DX0MrO0m1v0lIrkMMovcM3kGZCaV58Sak76zb5
NGgCHAwh8JuVlepOdSMpTGOw9i8f60tOUT6e2icCAvISZmWGfPWf6DFZzTaL
EWkPLliaoZuVMC8ANZhBv3nxCKixp+VCS0nrfQwVPD/KrJ8uN83N8R/apsrv
foJnToZNphy9MSPozCTUQ1fwcbo3+XGvEb9x/1wWbo2mVqm3OLR/9RVPPcc7
fDzIqVy8Y4DuwF41jqSVmpS2BRNF3bGSmLHsD4/6RFvhSZdwofuhf/OODuuo
uMfgrKm8Hzlq6MghIpBh3KJU8hOiGuJljpnSUemGXx/pAfxEjdWmx79fAVW/
dCySTF/j9PKrR+mSsjHATHAxGZzosUOr1wkPYZK0TTJlyaeO7ZjbB6U5VI6Q
y2kvkRH/4OSvQmXHBZJBLAWniupdfPMcN/Sfn0mZlavkBDdTOdlkMtcgR+yE
Xq1JzBx5sCpURLdWaZj+c47RBaPuqtAnIEy2xMm2I2FAXqxa1Msf9I6sRu2O
VHSJmRSSGG5Xb/+eEb5n0IqMR2oQBjjbGQ1UZJ581Le5mWdXYKl9Jz01bRxz
AG6c/s1s80ke3p3Zr31ISBWpAijVVDerSzVR2QRAuf3AvgjYIxw+H8ZH1mgG
RMEdNG9X1YdvIire5R6UlPjQS/yB4tRcoVX16EhL2e6gLTCdSKv5zhpajcsz
/i/zMT4+/xpLEvvVdufjrsO/PDB6LrUKzhrC6mSUOizgiExRA7lOPiumOT25
75dqEIuswcSUnSBcZW1onuLDFm7Z7YjrlKNkksrqrJhaI/HUK3gZbDb1/osM
azsH1eVDXOuTHV1m9RWknd1FORbIIOsTa+9qiaQFjI0pcO2Y+rJZiIN5mf1W
4Dvj0wzP63r+ulM4tZJ/n0ESZky893FlyVLShNEfr0pdnMmkOVvUeGuFa+K4
HL0gPzpzXzgyf4GkLRi1rvPMEFACufh7XNkyQWUr9eONkn8t0pjGx2+MjORw
EqNqs5xvFbJZJTDKlbZIFsrbsjv8tfmuOzl0G6ryeqXxdVHrVL2YieeVlRTT
DhzTwGdZej7adhp92elCLNhTQ9y7YrmaJszDj54KHfmtGdlFet/FDGcmmlfq
XQH7g2oYWDoOIkcOgjEzMQ9bs4kHMuLqsytJvXQzZLSNCR8b8khMtl74Za7M
isVupsHIIgHLQzkt6TH0F071oz6KwiynZjSpdfcjB5BVxmpXOtcEmyjatjLZ
rz1tu6i8OjCe6QAz+ggPslnzCI+8MhBdpOZVaEcNM/wtimwucubaBPSP7YzF
K+GFTskPadWnqEpOvAzrYDYfz1OKhroSBpetlCrM3GNFWp8IMViDd4+Zq969
w6l29N0ABKrYMpn9TQKAFrhNiYknAPNYkL+56eY16ZOu6NjOaBOIiZ7OGIQn
juhNSzV0HHs+URr3nbBREMNegh5dvY+nd+35t8hE887aX2oNsBF/Bt0Umohh
Ic4WVbhyDq+syRMlnpvxA4Z1VrN0PpCTue0osqaIvm3m7aKwdwUh8f50WolQ
B6LR4vOZ0VKSzGzm0Rvc3wM1GgJ2P+xoLrhUIselowllpWtQI1YqpsHvozqG
KYV+0rPW6Oh6a0d1itplobN61fvzwZOC5g1eK3ecz2N9X3ECnMYHFYZdz5yR
/HInmP3g23B2X3JLSi2xhHfAULuo1BBgVvfOn6xPH6H9B1/TxmzZW9aW6SV4
ucEn/EbcosWgcmvpxOlFJc3+JAzf6q7VqiuuQFIUT5wHPPCBRF0ddUpYHKcP
sWBomV/viUC4C0x+m3kduFONBxlON3ZDtvVDjCKUnKG3OBuWtZez3TuV7H8F
ZW9N3UXsU7iGRzHUraTgTZkfR5kqGALSrro0gNGFam/aH0Xg6gdSrXDVdLmE
sZo7gl/YPr+m1RTbJlmZaMZcTuvK+N7mV9MnKA2vyTAQ+6lwrKLTPK2PhgB9
jKz5p3a1OmrVV4byc93WUU4Dgc1bNQ2gSG73kZiEmYVofp8Ds66sZhrblnhR
wQR06MnncGiXdg+EMAzCyMmV97iLSoidGHaqjaCYN8I3h1wUe/cR+5LHCOWi
4pQFlpaEYTAdQsrbqtmEzR3/bHRR26wBRSangai0eYlm5A+u/aEadix6fUxr
SHqPq7TAu/o1O7+sGC6cOJ6ADLv4P2xAaxEsYpd5aEnhu9OqpGiijMgoZh1+
goRfziyj9NmX3GylekF3len6YQDjynF0KjOwXui3zzMgsRXGZC5XgVoh2ORa
IOLCtbz8WlaouROr2wGyV9MSt/jroVF/FtoVEYWYNg02BjXZiWPOCbKdVWHq
XbVReFLE+2a1DW8DSppyYXue/mC8GD+eiZYgc9x8dRIyl6HLDFFlwbes7oLp
CZeVIYVNCCYYQqvR6raT91/XHJnhwVRolSE7KbYK93q/x5FhGpUW7SWZq3Sb
AYoSKL3Dtc8tucOGSrd3JfpMclDtb3qbxYU4gtYu/6a+oDaUbPZ1+15k31nx
Rrn+/WeU0RMBQk4RXrnDhdH700MqSaY7Gv63qydbfD5k2wJweBxTLm5p2iSu
lQGmw9dmCT/zPfJ2iOwekWwbWOTIGd9cTAkweF7W8k32N7oD2SzCS+KDf6Zh
qFjvHfaRPoL69Ym/C8Q5BbXqLjLsFu6Zbpa2IiPgts1L9E6iJq9qQ3v4/GUE
SB8RYww57v153tYA+59ggmJB50KKUdujhjUMLjAYcB/I6vYSz0Ghbrsyd1x5
/tW9RZKgTOyVh+7WBTJ0gL4kaV/3BM/JLyVSR+ou59oYqApkUiYD8Da20y0j
WyFWxTf+1t9rx/qbSZwwyuzT2MxbO52HoVFHheyWfP0VbeZHa67Qp1NruAkw
q7Xd0t20mtjsv/51jvzS/pMClnl3XxMsB6sDyBvfjTzqmt3jMmClv/mfTl91
+m1hFBHAUHPbQYylL2zdE6+QRYxs9HJcVja0X9nSpI/N2O+v7rmvqCnutzU3
xvKqXs3w+GqjjYRd7/SXQcQ9vQg4dhIEWay5sFmOoVqpp89yqfhdigUiilxs
XSdd7C/lYYRCid2KC9BGd1Oeua6ZoJKSYUx1poOvXztUuraVuF6F97t20wFm
iLt9ErIfBLaTI8yhmsLfrxTgfdEvk/w8LIlVlq6gEv+EbI7T833i/UwJYBfS
HeatqgqZTTstjHaQq/hVKuusw982LnOGB/0qULy4zNFwli+K2j8UFySwMD2/
/kZnL9TEMPBPI5e65fzjM+KgYY9AivJkzg5hAfej7PanQvqqIFBHhhQfUrGk
5avqrxjvznn3O7gLSPEb73agAaM9Lp7FTUYch9NtVNuDY4vZRj8QnbsYmnd2
uFTY7ErtQTndDzV/D3+TBNLRKBT6Dq4eF6CkzeHUW8HTMMEo91Bwm5ZREjoJ
DNxzIWQuyzRYWv0SLPjD8uYUnylmLIBdignbJ0UbsVLAdmYA0ywlWqwbZAMA
CqD9IM9MJW6UEDKBfoJQG0yBU/jlTotEZAK0sUgQbL5yV4r86Y7OUvHimbjq
JXotHiNDtuVd13C4LZ2YlO1JDVF87iNadZzBPa6yzcI9KHBMBRcZBveHGnCy
DAlzyPVT1RPXhDfMLvq3VVHx/jQHLhQ17hFi6AJJ01SZhui1yBvQbZyKi8WJ
chY/m6ur1DPPQgkSRKpJOVKIhKf5lGsBDul3P0XUmIciOxTURH/OeEFRrHhh
yd3GAobp91pi0AKqJOWsY9HtbkwIiS2tWJ1huYlGvQ6Zs4HBh0t9auNFAEcb
kqUPu3wlOZ04PyLhTjOmXfmGVW4JXsN5AiF1o1X5gWnEmAg5QKMIfhahTYNi
RYR2cPBhXoEHBOFZx/ofnUOK7h4IXKKjyhsneB35tmyayRkOeN5uf+89PJLn
tLwE2HyNY4SMvnijZ2ngO5p1CXOlHFZB3TAdvjA6PDXNCzjCzc62CIUNy7P8
4lPPL2efASUMnfqpB8PYT6P9aUteQKntt7pWdaZu79/jGVBpXHwTNxsKsPK5
y7cG8nL3hLnR9mQqMRpGtwKsjFFIfwak18uLNfrIlHTllP94Btif0k58iH/Y
0aZI8s95RLXdbKUGdEO3omhAGCHUdKbJY4klCd0bdmgK9zm5kIgRUJk/fW58
sU8LTQBVKJWPm4ModwkqS2YKEuUerw1KvYpKdWizyBEiSWfun9MM1PxkTfDd
TcV/Yxrg3Ekbt0JsqZA7pg+M368iocAUtoB5LYD8jnjxsAs8pwmj7Hbs457x
z4a//Sop3RDo6uU0AgG7SxMza1Th/Wo+2Azyq2Yq39Al8Vgh27AOq3RvCBY8
2h4WYvN96i0vIT1AfLmNssLUTgE56buQMXwJ5r2PwAD1D+Rxy5ndB2IDg6xU
bA/gi997e9h6CWs77oiM2agMtHshAIgyfSJZEnILNWa8xJR70MLGgLsfJm7C
u8fJf8bQxO33ZGywWfqoXCwXlJoRFleGYelcQ0rI0IQlKzMuxHDjg+m2hIlu
4+CclysYZSGkCqaxWMxTr2KGv78VmacONsFP3PWPGyKmOfIVgxSqjAKa8wx0
aaG3ORE0cNByVzkt4Oh5rlBEObP/eCVsvqQpAfuivGL3z5mL54FEtXkF+7/v
d34mzf1KE8Oo9UUzRxcDzS8HJxZ6oRXW8OnZZep1h7Bt/9MAYKdLotuZAcMH
rKOD376XkylxSjPRb/IdzjjNdQVU74WQGIW0PabX8pr3J2QtOw/yd8OUmOYC
4s3rfcxqMnTJUJPjMALSftOUWusGqkMWnDaPKmnTRTo4WB/B4ote75P1LGPP
KBW/M49oCI9j5PN66loiXWV09WWACn7msT270id8PZtBs6laiB0trfdW43Hz
0a6BFxx7bKoSBSXl1zdYgb+BefnmGt7GbcPPhasNSDoWnTGUiEHe8sr+wad7
INdUIT+EeWCf1PADK50N0xqPSKuRFuGtRfwPzR4k5kVEtE41uAOnApKSKI2R
KNOvJP6osrNbgoYDIUKZLGSqM7cnydU+cC+Ft+KB8fbBqzuvwbEBShA5/eKr
hwj96TT3yGDWNCgmttA4M1L/HQfXi5BJ+kwTf57gIxDDWWd2eyWMNqeH8WEH
jTaQQPw5tQLDRVoMNtFiZ1S8D2tD9EE5RfDZcP8qa+5+Cus6k0SHFr4UzylN
ricRy5j1DGijPYYWWssBXG/jLMz//bZa7kUoEHdvXHLQiJhI9RvoXykQ7bnv
cjWSlsQYnf/MdzWVAq/UfM+xYe36pGpMDi9/Rxg6Qf4wJTVdwLqIAAY1qbaE
MN78PzHRAuR+GU2e70+HGnxLrDnRkpBIovYOs+HFcUFeV7uCyogwefOt+7FX
kHyFTdY5jwOKtzRnElw58eQbhyT0cO2kRoSOw54/JNh8wkycfUO4CfaJdFBk
L0iVERS9fU7+hsE43sDDBb4ldj20q3Se2cuCo9yGU0zKIjeOt6fYXMQhSHys
kMXgKcLIa3wo41aTP/FJVlONNf58qpykagbW41RLJQIFsuwyLcbMctFEx72F
pvZLx+Rn/LQy50H6IKCmYwBYnyqBaDgaggTQzsPEiZz943NFMM8pKBfHXhnk
NntbOWZQ3rhHe/Bb8FWkeQBr2L6OIS6vb5e8Zub9ySEprQYBnp9Ha9UqX2KF
JPNHw/jXZbFcy+3uKMimyF9s/2uiD1I1YBiDp1Ll30UGCUtAe8v34zT8XeBL
dG3v7sDUlBQBT5tz+yd+U5Q2Vw3HTfKfjHeuT1JdbMO08ZCziHwXma5Lldh2
ck2UIMhpI5gBxdJDfzHonGytAGQ7jA2kzuc6D7PyZoiqsa2i60eTFYc3p/vI
k/4rMxibVJ3b32yP1lO855C3UtWKKQA6dySC+fZRfqzEQAlz6DFHydynP0lx
y7BA/KfA+PNTTsMlfE3pC7HW6UXWDfwrogat9Lj08/+jXtMpunqXexOLVEtW
LwZB8bCnlIGqQbozUjfTzphgw79CXrmnyxkhL2QlJQBcxNSxpYspF/mNyDJw
afzQFpnJ3Cy1qYSth9frcvWA4f3i5IN/rbi/qpR/syKsXO8b6AeqZ/o1MHAa
jhreYzxi0UCAeZwFfcitBxOGrvfJxQqPYyt95sM/6jUuzeoyn9A7I2hi0VZb
A85BAJU4v+wBqLOgfinC3ou5NxgZCZx5DDk3M8FrOT8Q1ukTVEL3Ht+QcgPh
yqHsJMLJMyAhdsYp4XtblOIxscRSuDXCEcLA1b2VRjSTTIDkUBxpixFw14j5
Ww4zJKj6LLkIHaZ8IH5imhNv0JQ6asBI6203SIH9oZ3dsBmLI5ownlH7fhkB
2tCoaRE2/JVuzHkdujtZk9C6hEHkTLOEVBsQOooUEOt9pybmnHrITYs56GTA
ab52seFq6jz8EQONy9FPVyA7QXwiZgIfwLyxUAz5MhDVqlaisnsdn2qEWtt2
ylWO15+7o+7UJ9LLSgzWLi8aLdu9+7UbSrbmhhAm9zPEx3B+r98idbdu8fJ3
gAOADokTk8k3UJjwtS/9p8r0RhHKQYAJc2gUGhwwseQk7IrHTGX7IBNRuy1o
eydillqjLB1IequCl0O0bHxh0OXX8Yti7+doXWJTGmtVJ6JjgcPOwtt2E34h
NMOu81RJMv24wVw2KjfIudwTgbfusOy5pTZGyYnuc9N6Y+Q3XLlMZLu+nka4
MV92c8IQOixohLfzxddzp6awc0mIGPO+mK7cCj1UIoVTBAt4s+eNG+vrkMC9
OaBf6Ehwliyf+zm7gq396enSTmx0IAgjKJ4Yp+qJi6oad/rh1wBDOK8d7unc
QuE8NflTax9R50mF5AQ1Ds/hT9sZfThNd1p3GKvYUWz3ed9sa5e68Pa91H5g
w5m1v28p8Ay0waj+Y+4ppdlhiOlBAidqwAZbVQbnbDW07CR0nHB9VIw4bH8M
2xx2akTf4bf9wxbqAmzzpnvf2EJ4AstR3+gn9NHam71DGgJFxjiHSvxsXC+J
J+jStv9NgLrRimjm+T3LnO7pJ1jdZjVS2KQiu4ll/Qwq48BTbfaDO7dRv3f/
7UfrZYZP4WOpcjl9VsgPv3cvekqjOO7keKgq6FFAaArY1+jcqjj8P7ClWD3e
MjT4MOmKw0EFxb6yyhP1e5SJEw4H9n9k0iJkuZrWmfkhaRW05cJLTH6i0Bk7
U3w/TZNH/pwh5XMO1wVPzOKqk3ouD00t792QJkd3glxkNowklFr9o8n39s5T
A3IUUBALFtZLwvWuKWTNdlD7N7SvkiH2z89dliuql7JblS4E8VxfeYjQVeWy
uUPbty54TrZj5N7aL9t43jaJ2LDkM8cRnUETJzfiLdBH5esN6ipHImeWaSWU
P0/qRyrwNkE66fSWFqruYArtJ4oGfvNfCE9UVwc9l1Tc2OujuKELHRd3yxlq
mhjJZllQXkhcGzhNX9T1Kq17MKp+G0+0YjEtAwhB8DR+kajxpiG0RgxXYI+W
X3/RVEgm0MdFixU7TXyU6qyieoHK4mnMDwGGtlp3u8gQ7TiK4pX2sgDwoxKh
yLDVg54z0XJttUFgyBhQLjJ9KDADo369yprOsQ4ljvukg8ydMBx0u0+U5uHf
5QZI8f8UMtszLUcr1VMu7McHtclor+p8NDe2ONrSdtsBIYjQSQS9gIQxYgkF
yoJVhrBkAElXXd3TJoEn+O7tWd1lLpVrtZH2+UFIgLhpjwFnxKATJfm37fso
LXG+zEUylBGNAFdUMV9gx/Ul7oPHuUJaaHKeFSI8NHDB0tX7EKM7FHrF+fuH
nPNaUVoKQ1Azt0bP5aeC2zd0cF9skrPnPTuyelVwkviigApSCdbhRL7bOOZ6
7IaDt4SPQDS4BvTEYDesh/I0F6LrJBlQhiL6VwCMjnnW6HjEDrbarbZMiDAz
58X2cGCEa7r9gRg1lE1EsHEOqL739uTJ+lugL+pWdGJzw5mZ+WRj/TiqCVoj
q2poeqGzA0qfawloRBs9iBh+9qTFI8zT/Rk3rJrBOMqCkeCtsCEA8/7z6kOG
YUyIoAkCL+LuiiQzLNGCQ7Fsd0rpMIXN5NW7chEesTxKlQ1BU2O37Uaa1LPG
24Bpbol7q8BJbinGvJrzYC7j7yhArf2kKJXnHoMx0VZ8nWcM3V+XqsBOM0er
61tNADu4mER29K7EcUKgWDJOr+qOUQPTzlZFEbqPTTDUSHGpDinUP/epfUp8
+sZlwzdfo4gYmjEzzUWY4yeuumKJzQf8f1yoxz6PLepwWjl0a9oX/0iKUVa9
PmbQSHzuHDgOCpFyb9NMg3UvBFOWHKKeKqOOrnLfS+l813JI9mDOh+wLNPio
OJPnMavZPJzQG5+ca8ltnz1En2yOk3PyB/tUKb1rVNeoRX7O+vYSx5F6zaJg
jp75pQkIGiud3eMoGddozZm4Ohf0ekuP5GLBq0YkwF/B8OOvBeLq4SwD62Ou
Ac6hv+W58MZxXy70xZYDUPjuZk3wiK27qg4TIA9TrK6kxjM92JlFw46LnDHW
O+iQjSS3LesRPMbfz+TbMsVJFYTQ0eDLLF9J5r6/pGMfKlYYQdS3B3JxgxOA
yDE3mWQqqfUeqHSyt0iJ4NiIqbMWBcycana9VfF0cChOd2zWA9lfT2xhiuEW
3KhEUSYGpOXd76Hejlg+UAHsTU78mBBaw/4WOgzFvRnP7S0HNX6Fe27wsS32
qStE5C2zHgBJSXUKWNEhnnrc9eq2VEXo/vB/JwohY+Md5ILDulUT1rvjRoqL
BuaOr5UFZ/g+DjFUePCPPGZiLaOE+hLxoATXSLvaf/aFnWmuZwRT82jcSRWs
TKLRYFUrw/7TfZHqN36na0gIEt6awbVLwKIS+/V6nFjYfStvUCiZw7jv9zxV
p0T/BU/QQX6hFE59Z9UmoMIQsoZPKsYayJ5MHyoeamkL0YqcoXRJBLYky/5v
R5Ki2NEv1yN8OLJ6A7qVCz3fTTT7Q9karnHj4lfVEJgVjuA8V0WOgxVLtuxH
jOhPNga71P5zYI/PirkN+Cuyq1dDQeH8txUjHTJb1a2dmMAQTk7HqqmPeznV
58DGVDiNJh7jwPppyopPG7PBJwuJWWoua1E6ex5ODAb/65+Ritw20a66l2Pk
aTzT8CRBdAnkF5aaz7UrXw6cxzLzuv8/DKxPrRaGgbJe76oIA5PRvDjDGhcl
7oUNeFWrwsYT8S7p0iwKKmYKjZ3iEdiPcXGlYwPM/B6HagMZSWmGNcACfsAI
4fUGb1Ur9O/KVDj1cJAwDTIqCFa/2wKzKQViqwOPLdlwMrKtcnDUXP0MAcBd
skxToMIAekQE2yyOjHcrLFGKOWN9HDgeGQZj414fxfPa679u5eLJv1ZE4xve
0U/Ks2yDX8sW/q9oNBv7NWOM+373AlmqyTPo4nYiiL8w5cnWWeEH5s2bVTKY
kRd4NBJK5fkVzo2c0l8iReDrqlSZY+zQX/n4XfhnxpfmOZEAFV82R/+2CwDd
nanv+M0ufnjbcYYOjucwhiCHCWCg4Mh9UxHIoCKmJugqSAI5OTkP/27Kni+W
zE7yFUc8Fy610ySoCDlqEV4fDHhZMPmWKYX7YPZO+UmNSVkhZvYvDSZP7gYu
8FvzLjOIOTVk53kcgIj6dZA50HBmUNRbA7c21Lf5p0AMGCD/ItDrqSbndx5w
pkPcvgk8u3xmz0+F1ttrGvGGWaG2Ch151D8g9zWV6H99rZ6SW1CqwffyTJNw
Jq6gt47twY6ObSZlhGSJqmwxS53xNkqCJhRILY1ezOmMw/VgH571MU/vEjLZ
vgZbUS4Qdcy5UVy/vrep1bwo0Wy3fAXkeyNk3upicBqt0NaOb/N7aCLHKqUe
BYCN1G/6PvZ67AP6P4EdfDQJbhfq1qMtJT8VglTq+iEQl/Y/L9bdsCVciKGX
prydIpWJ3At7SmNYFT+AN8g5Cqs/ks3WqhxhElFXOFihkWRbAc5LFuvap7L/
HwTmM5R8t5z6syMQ+MCwdCoUwmZJzUfSSlVgKUpM7NkDf11FwAGP8b/y+gyO
WkLdRsctYnPSn4PEvqveAP8lMm8TJjdEcvT6/ou45FKKGolIFeaZhCTrFaHa
0C8dYxKF6KrzG1UkLl+/Tv0O0ub/9ZB1Q1nJQ0W4fp22YaB45p1RMc5QacFZ
O2FpEotrR0j+t55HlkecT3H2sSVLrAOMIlfMaRP3ZdGCp56Q7xdegRobYELB
GHgT5S/eqlITMRCGe1Lj8PMGDdOMsNkQsYAWKkUwJpfC89cyYhyEDHTEnHyo
t+MqjAdtwusUPnsVxpeaAQQeMx0AV8pWIHnVpfr/9ZIw19l+shmj+MiYptaw
25BWg7CBCqdFnKpPE5kH+Ml+nxg/W4MTh5DeQZvu30rDI41ExAwWIgKAVWqy
/ywpHbEY2sV9uOo7o062w9TBaHmVm05DWd+Vsq4EdTNye2OYZvguBuIVEy9A
cux7ibXnCuorq8yFGZX7Lmm8ivr3ap/aTf462pqC4bngqsg4Km7jDQRV6O9a
K8t7oddEu/NJ8JgIahW28aVWNPXm62KJaIczJfM7TQi8nQIOLm9j87X0b5DF
yrWckCHUe0tkAwlxDvQcUllXiyIcAENXmstESDbB6+LC2DqS4fmxtCeuaV7n
gm2JO2Dy42CJVsI0sL7GMAdu61poBlN1Pjp78EXoaeNczQStb1LIR9inBwXT
cO3/iBB7zWt8qJPUJ5zvp0WayaG1dmXXR+3XyXEZ4HQ19uxOazkSFd1DmQwq
zfZ0rqch6xVPXab96qhkzEIpnzVXIkNV8LtqfU2EavYh+BTnDYu7dOjnmWe8
13SHT47u3RDj5lyjdE/esydrckYljJmv6aLFEOdkPkgHCUoxZSKMbgYDWIJd
Sq4U/BslQFloM1F6/wkVVadZeAWm59YToPN519EijaDLsuZXW59ILfiNvwd5
kqzTq6puSnfi6OJzbAMFKYM+zvK9kO16YgmsbXr7/OM8EYX6o9nESy/ek3Zr
YLb/LLbZ3kbO0toex//tyMz2EoDKVDB7Pa/qWjg3pClCUrVMK4A1fMkljlhw
SOBKUIYZ/qmu+8pVIxzjqW6G7OfOS61qMmhuJmCTpNaPGZ45tOXgpJidUrhB
UP3xlSagCWrlY41pWG2bUUQBmSwxf3eREekCaPcsXPjQy7wiTvRBRsfc2Nrq
KxT6pIIbZFR9F02kfNHgJw/aNUeXN5YUHm8Mi1bhACuYt1xETBNfDa+Tqp4q
qf7gysB84noqoI8PPxK2kRgFKvirAAu8Y+obNUdON0qmZwqSZ9zYJ/J+AyEj
S573caGNS+fhgO6x8/yBCLxL8kVZV5vSeOCJPCL9YAHwH8ue6OZy7emXcucq
q1fX9bYOI4o3rxSiZiRpIcvguQ7PsXwDatBshMuhuhyLKo8LKg1CT/No6RBa
bUqhq43nM1vMgF4mEqqu9iEWpUvbtZ8MVXECg6MH3cLFHHhLMFfctr5RRNI6
GF417CX5bMRyoPQpkh1ulhsrjknJllDwR1DT9hoymbBMM7ZEH84nmWIA2pKU
FyzfHgcfD321f7fYCDGWvNfcPwRr/xl0c/8MpKIlg+CEQrjrY4QIBXUJQ8Bf
JNr8Or4vQvsledHWrLBDpgnxqOvrVsNxdl3S7ZhApRWNbDhd3kK2vEymZy4n
MnIH3iQrGK4v7GZriXMCmjGWh0KKHOF6b7Apn0Az8swvIVHPM2IDKWZU7vnU
eOkLif0BcAsd72EvyaglJ4ZKA1RwQWbpMhBJDiWscpBuO7AhR9hL9kqjIFwU
knyJRs3oL085DR/tor7aKhQtBpTJ/OpH8u7VJNs9A4EV9bfIjCpgqqf4xm6u
UxblmEaZwDl5IOVul45it6BZDI3ns937fVXLk5BFWOJuEJjZEf1oC6FM5XK9
cd9vhzCXIDcsAvSp17vuweHdGwApoDMw339ycWzLAYFMrLZ8tjW/KttFUYWw
GQx+WC65csTEbAFtwUhQkgCKtHQyC4LNNwdQQ/xQaT+CN5OZrJOyh03OQD7J
23TVqbggydUB1NaTDH3dc0rgEtreJg0vRDDOCBTBeeFG6hle6RRZSkPQXikA
x34rENyqd5hyHP712izyeFej5FxpjsIJRrECt1GTfZaUzcEfGXcVwNRWeTs8
vNHiJBA9tpyvmWZLZx9SDvvaVf7OpZj9eq1znA09WLGrwi6wQl740i64Vi57
26Frx6slpbYFa13DVEpj7JitgtN65a3VKnO21PLgS3W8c4qz4iJh+5dYYolY
6ycmbBCElBiFq4yTsVyLpRrEHLpS5lJerZPj2Xs4GlL39f8YVoR92Y5GapGq
X8mOtmeR807HEyQehL5YjCVNeHVtqIqqxS4K2NXnPbwwrSHpqg0/YgzpmFwt
SzocXTYciTq1gxiLxsU8C0dJCdWEdVklDIkcG8J6dWU1r2jbiVygKmce4PkD
KpmHbmo3u5jT1oJIiug5y1okUJ9N/t4dsL8+6hlMIRjRhKbvP8Pv8HzrOk8O
MUg/i9c0f4hE8xJM6meVVkOVe1FYUzkSCOr7mMHDK67repe3CmykC6bF5DEX
JfdELCqKRsRHLOrw2lzUYyKqaTwIwiga/2RMydXGh5tDHHkHdbicW2ZwIzmM
9aA802pqCgpoSH7EMWRdVgkgNCGHDInaOMtjrGrlJGcG5uq7PjWwMvPSfRXv
1XViHKFeh+DMug4ofMCtHLy+UQ/QY6jhF47KDRA6NzwSU4d0ZjD9a+2ArUIF
vrUCzTKsoakol/RFAHRNIzNZCB8X6oAkyOpu72pNtVkwUhMduMKvLZw6cKAn
AAHJqQrrdpmKHBlIvd3lovpfLJx/jlVFoz4Cra/6r9P6st8lOc/tLDBenZLF
R1GKBeWt6gi36PezEh56pMi/Gw8VKxtdt4FWckdx07qOcPHyqm7bLFCQaQgF
wljUGpiHlJQs9q7Jux9TW3oF03JVAlDf7yps5dGsP2g7ODc2z/lIjnO4Od9Z
zBZSgX/nh7o5TfYtpAW8nCbJB0lT9ycTbNPCrn7ulU1d/JX+AiWoD3PWgeNs
J43lIiiXoyq6v4Zd81cYG9AMDbHRzcfPi/Rag7tUe4WcrOCjMQglHO6eKfLN
8O7Ld9pV2PlBSax3mAvwTCiDrl/u5SNBMGf6eRLS7rBIrVLbZIByp10fyoJ6
d6O5qdRT4WzbkFCbjtKUub41gm2quToUQJxt9RjlaozHFRXFIYnEuE42ljgc
HcXMPNs2G5xRHyggx/gewP2s3pAOCrKXgYHFO+WusnkRE6EoOjGFVUr9SgTu
LMkltWCg9Gfbumu+NrHr3YxFC2RqOLgcfNSVvFpunGE0IGiOasNdyQkR8NxG
YqK1BZ0WuOx+q2Prtbi+RDXoL7HSbkVRi6uW19rCgUGXWA54c/D7/k5GHEvX
XvSfzKR5QmwlKLUk46ZBKeE/bWJuge0otacybTLOuiuX+WM7hgjw/eMklIMe
Hl2vEoQsg9WsLMmwEXlAGQVBq2SQ27P6bBONpUCN2OEy2v1Yuut08prYH7zu
Q0EMhBqlEEFEb2ZkI1bEJUGgEDjyNqgRwswyV9kTllKtifb87iwEc+UmCh61
vqug/Hj02+45PpbzZpzu+BqL86/yvwic3UbTB/7vMwnmQT2J/qR8RsibaV3W
eCOJzMIYYbfmwhHfPLYFMS9jaZGoW/pSJy3GaOmqAFx1biVbq5I/2o78cofC
O4NtFI32mF9ZygwXBdrU3D58G3mRuEEvnc2mgIMs9L2ftS6P6Xei0wLwqySp
rv2/2VkQqHKDTz6DsrsUKMz80H24rG65ZSNapsm8uD7j9Buqqnqly+bDjQnX
B5xWx7I7l4MU/F3xHs5MEVl43+QjUB32P7V+QwLGsEFnIVMYgE+do8YlNLgh
ZfXlNdRuC0qiS8yWT/h/tUzoimZmeX8Ox6tDzM/XB7skiGboDtRyE7bur3oT
E7lzA783BIM0UixuAF6CKxzdWmudv9qML3vbVcl9XVWxh1klrQL3krv3xoXF
3H1xUB801DpoFtbkp4XKwNa6INr6y651aixANwogSLOA08ztSILCsDf4G9e3
qgFGlb49lTw5ojvqwdFIpQxDDPGgv0KccMMjvaBV1shDag/oGlxAd0sA7IQO
FWNoNpLnWUFiFueVC+1R/9mt95S9L5bnz+j2R9ZF49CoEjEanR6i4Pv9+wVp
50Amn7V6GvhQn/zYNkVMxWYHYU48dG3KFGOtOrbJhbYwvnr2/P9nfducyktN
R7vM+0DDoSpOqbTVe2Uv26WI8p96aRYJxI3bljTEzVPwiyo9eBMwKTdMjz0P
ipGJdTEoce08qGDAZLeSHqiCjZVf3iQi7w2U3zlrN16Ct0Dxfz+PcAOCf/Lo
X+sAyenAzier8QFNDFujEJ1uoxA/+pfB5x4qc08nZJP2bHSM2Ccx9tImwnlB
yrpUDEcdWzQ5MYCac99gLttz2UzxXkOCyFGS2U4MMLucErN53LJwja5rXGjO
OgEF+LE1soW0I6YzT8KjGF/XZ6gKxCJzZzuv4v43nDpqqASr+tAodWf4DdvV
zw/8uJWeS9zb0CbZXxkkNsBIEBkAfxGgIAQbBMuPINPbi5Q4S84KBrFNb1d5
WlE5yfBMGJ7W7ADobcnbQrrQszskov6tDWM7KFjKza+swxsdXG9ussRpbAeL
vE6RZ0KbXDs34ME6/oncEc+9sPmXYoszWav3qA58WbM/w9kCfvDdMakiEQ8c
O3VFAuSEeSFa9DJ2EPd2d5q8FdhhPevVakvm/p/9Pzv4n5zgslyrNZhlZEuk
VdFzNP9tNZgQS07a8MDiFUYDWMoUu4mLNtrRqQ0sVuNWLJOmd6H8WfRMMgdQ
5cbhPamsmL14HxAvgz+rmKIA4u0bYeH7tkw4uwr8SDhgqxlhc2+ftzuNARGW
EX6aHLvv9hSsajBB63EJiCkYvevoYbVRQqs8Fd6SiqdetmWa+4k8VxXeAMWN
1O3H020i6GCT200IEmHW4BkcK21hX5ND25NH+P0Gjrf0yZ2MO1HNQ9DHcoWy
NJGaXzST5iW5lX5TUWY/rX3atPk47TO8nMfSjXl/Zyn+LoGE52EoKGnSJ0EH
zhFreovBGUz9m2Y0N2npVpC0PVWMcqYwg1Lr/f/YNpim5t70h37ky7HbuDI6
K49rSXAnJ2BMjt/63fKsOn1SIDuNKzRjmQbTRqzZv3zgUF3eBE3UU4sfdoaw
vVUDvnsQKRK0Ji1fs1R9n1eCJNM2vGwcMbumSLPBdpfOu95NjvWfw3BOuaU7
mulSPkgyYuEYV2uqNDDLqRw6rCoMXtzvcwPgAfpdwZfP7xGdquwaUTq1llg+
sZFKV5P2HWpm0t1b5wZSeN1mUCaJ4J1yfsNQt9TnU07GuiibxnXPY3gK68HN
sN8yWD6KaTKceOOn/6AK1PKFqUbMxRVOgriH4cHTN5AbebFJISBDzfPPWDzY
JL/mhihaasyb0Mv1MFX6AxqQdTscsWgVpz6eJ7cAZ6aCb4g7ZuBm15D21nHk
GRkHEfCuPRa3+WbJWeJHBx8nhd6a2oFPjws0WCC4D9D/XTVJTIxcybzxeFi8
AMunoxxEtlG5fWNeuwhXeJBXNJgfnrcMAccG1bP8jg+v0bFz60lT+jRTOc/T
6OaBvcRjqGF6bSPhzIptkFlWnS8M8an1szyDUrFY1/jSxfFMfK6TDSi0nvEv
LLHCt1TZjchMUSwW+JVdsTFIaG8aAypUbw9CeO8oppiGA57sIJq0pI30vHuE
u3X18O+sPUhdMjI9RE4AOOdL54/kIYw7MxjaPISNUwwIMr73wYJBB0DjqFur
NQbJVwedAAEGgSpCM918nNNHbVoHNeWrDMcBsTcCSGmvkoFht+CWJQmSLg67
+EqR52C6mCcqf7clX9TiqrUdx6Jdv2XbGvzwfizhK+coOdUWVzQ1XV2aFPtl
gFwkE5N1PHziSsckDdN5PoHmH8uPGHG39SJx+9vRgRTr/40LkauXjSj0pGEl
GLJZANUKZmdDrPvtCsmtzV+VVo/JeO0AT265/WGw74ySGJ9WsBOcfUjR62rr
lxnl8LtmPGQRgrCLA8NyEuBoMnirCCz89xs2zzBUPTtQUjsGPphJA8ei1t4t
5yHLKRRkhr+rxQ2qIIrLYBdi72zFO27XYWgB25M4zS23a/YUA85/KArHmuPY
LOR8wez+wS9r81MVqp+z2MirZldvysfXTosUwqE1wZHKh8XW19NiMt4mYtBL
pokvM/Qif3bVHvpg1QsyCUx0+7QdXUGYFU1bn6VQOFxo9qUU2GdPi2B0vdOP
szJN+qbA99hwC0gKtx40p3r9PTo1ewK6K/pUIRzvxzJ/eNXk6qe+FFLIauVQ
hE2t3K6Z1Eff1hVPH+4wbBe9OEGoegJL5XmIbsLllx/Tu7gKAOwH5873aHQJ
nruu8qY8Lt4my42YzfHjdOD7NAjy6PLM0rB7hzhDJ652MyGHdebqhrHmwksE
F5dLmYvGzAXW8xtsGt3+Bz7EB1x5db8jfOi1YEVKfoteCureck90+vWxi64s
Gv1EfERhb1PtXjcb0KCqBbwyaGZsEdiZpWwL9sy6ACo8zhJ1mfKpkWFh9Dn5
N/AhaRKyA8/eJZEpybj5EZuMUQ5tMfIouSUJNevPqk2rIRyWUyVTduyxlpV/
34OARk4R2/GtQ623VV1NE1QfTHi+aRw7IEDMP3P5PDc9EpMjGTUoVcQ+WL3f
r7kS7wPBiVkzfX5x1GFzAO3FmCwaokoFekPHjbeejYLoU63zT4QkVP3CYTQG
o1y/2j06BdaqHOErX2cndYJ/gfDdMkEyDSN9INYKCGuGVAQlBy7R6+wOYYHa
6p+OJvsP9bgjuzhqM9HPBAB2bAGUKhV7CMWu9ivbAMLCv2JgOnAUMtJuCaJb
ZDvKDfQFJIAeDxlwMtfFl7y740I6D8yVDGT8XdkeOV2ljH1MeQtqhvafM0mS
a82ydkcuqJ57o4SLa7ey5854FHIoiub+ee2mfCvjIZXeGm0xMHR8ynmHd9VG
8T7OaDi+P26xKlGgdhlsCD1tC67MWz6mScBIp42+TbPtZackL3YJRW7SrKVU
rg3pXrKwl2TSE2B6VohelqGA/oY9wsInC+V1GO7pFtLf4QFTrfk9a9z9HGIk
sMMrqGDaLQCOEgv6ehCBqic8QEoJ6WvZAp1jWPjFwP4vvor75mTJurjdwqJM
7qBRy/BrN1soDyqWqQ9+nomzthvMYsfYN1TlE+JYdedWQqR4/el5MqGDhARR
4L7pexjbqWvAfj/A4HnEySknzPYF5ZdAXUuR2JyabxQAeP3DWV3LieDY1eEC
xuCFpDGsu8i9k5uQVMpHDsXWGPHnTtHLAX+/O2BGFkyoyn7MquB4weOtAAOD
TVoM7ZyBX+QrNzf/h22aZdpDul6hxCYgXKnYRxVVevUyXyPoYn/Wz6YthwOY
IV59sRyNoR1sm/M4ckqR/ejrX+HwDOoOXXX6lV0zrHtwb1YbQ+G5Md/RleO3
osCpj1Ji3iB0ni1ukE3vsSVXg84HwCPL6FclIyvNuz3y5VzygnaZFkcdwqGz
XnBxpehhxCI8R+khLXlMUCYFgza9OdrR/Kh3vaqZp8z4stuV3Xmg3ONHupO6
KPV5qQ8Io6AXZ1Hjhhsla5mTw9Gpj3ZLQBFwiHpcrRTF1GUT1titqg01TZQf
LDjBSfJW5fqPyJRvGxde1ORa7mo9wthB2KX9LDmRJU03U+qGrmIUWxRCuX/C
1r4Zmy7jdaw9MZ6IklEXCQZ45ox7ubqMSyO+PBg5Xje70N1b0us+Qx7vJSpV
rBjDSPSDvC4EtdX+CstdbZFiCJ0cJ83F07dHBfl1fngVqQKftNPjwH1Ni7Tc
i7qpKfCUr0N1I5LV0y0gV0cYJ2sdI8v2/UcaNfmAyFS73vpyugilpo1xy3yw
qfEuCjM4QFBWdBMupKyfepf/ve72N6M+rQi7omu//nF3velMilviKFalh3D3
ahkXiLAvsIKli4F2Iev3JaNummvACQsWriEDQGVnj9pqhJCEzhkgQYQ8rsZ2
ipysiYDhiD1auN2hdW+BneYfRx3BF0FPrQzbxbgNfsgp4uvkCpk5ki8+OKad
oaMCW0VEnxE3VuB12O9UlPXmq2ALgMoTu2PWleNSJt8mPaMsW8s7Wp9rU/y+
0ZzrovguG8cB4DPXmbzZauvEJ7h4XvrmaR1bZiFESYgq+1qby5RWo/93n2ah
wyhX+BtRGI4B3XaUARPJUcAa9UsTyeRkl/7e0tUVluZ7tyQo4iXCTJjMwZB5
SzKNefMHZ/8e2Nn2RbtS0uHi7mr9lOKXstRNoVoDnV6LvNnkq4U9Nu0F1XMi
D9oTlw36PiU9/Cph+PDGifqJ/nlb9P6QeuQEa9VQqa4yjQAN2DDtKl4619jU
9+3acmfnB6+XWmMnPaLeV35PuykejA1BBk2kpqjNJYiNBr4gJ35ZRWRt6gBG
WPCyAyPwtLNoCyTa2/20BkO3Y1W+4w2Gkgbpy/EYJNXAIDNY81oX2MaFOP/3
qc23ZvpVOZbaSvYbhmjMqeFZ3aQCkxhHV8eJqk/2DxLmDd9AnBqf6bKEwzMJ
PYE9gwGYs/RjsZgoCd7amvaQzRJ7S1wUZabxCeEMzGg134m8Xxoz2HBxh6nR
zvHBcQsAbR3H030wehKKUuPd3nJNi5M06fTIMBdgOQFP0fVdTFhE60OQKZPv
Eig6YhQpsbySFKZZvq8jv1OMOGdWKzeqAzLBWwPytMd0JSuSBwg647BmCmUp
6mLExRosOIDwrBTnI8lBkNWugMO0CeN9a4/aFsmwzmfAD2djMncuqiqp8LiE
g21mOUDKWMRbOTwZsM7wHDN4QU94yA0ybX4NilRL6LSDVQZcBO9Abo6SCbOI
2/gVEuR7kG2vVr7kFKAntTHRewFvoryCFPz+mbmvmljB6ZVhbNQ3rsarKiTb
oRrC18Kz0pdaGNg3zgzE68DuIkfTW5tRdxESFyUO1LAaO0SDFc/SLyAb4R1q
4/WG4niSn2oFQcFzxt8lwKbRgZfBpymxuDyACpFa/qGCpypMlDDsD+bRkrLS
sUiy8ICWcLnU+mrprDbzLk4XvdoJg8pKctF9nDQbqeSaTq7fIR7s8GGvP9Bs
uLO9SPHGSRqVVCpPwdmxsGx+xNFD/6wHfztPXGkygsVwsbdXJ0xN47B3PiFu
FGYfhkhM8aFpetpR8+rdkgNrHMUxnHpRZyxUWoCM3WLsKxGIvm10fI5kJKf9
6Tp+bOGF2QEicoPCA4ognRg2L71WD59PfNR744IZYQi94dzbcC43dkEzwJE7
KKFZz9xpvvHKGGDfbqzM9YYioj02HMWDxTAiileIOYu7ZEskUYLRgYaC9sTc
CE8benL71YMc1lDvO1Fl9S8k4U9OckJIxvRZXQJmhxpFmySgwbYQGyUIVj2A
O6G8jyMo3vHHK2006iZ8oEKzy/ti6DDJ8TjSXfAUyN7QK2TXebWxLtqo+Ium
OWlMwgtYUCkwd+vID4u8IFKSEHFt4kk6Lnl7Yc7247YBLl8vmY7Zzbq4eHL0
i/BmkQFyXQoLVpjzK+kczzIh9CfpXl59POhUFHn1wos9V9a/42v2o/s7UYjv
Abzj5nNy+cvDmkiGXU8DUyuVMUlcnyRVQh99ZJQCMzb29HOHuuuIqxnlFEKY
lWJEIC8nzjCAx09+L4A7Lavqq/tzys9xdXl7FUB5IYFpFI2CAhxxrP7q3Cj5
BoIYeooJQzJA8abQ1+pxE+pBg9QIXBcyUvEZUnSTGhMLnO22iIOI75fxzvkV
ISUw5bdAJ+RHFm8VW2wuvY2NzZCrO69mfro4uQ8lrzCTZqI2wNkGBfJ3ioJT
CvG5wOAjrVHYulxmhjx+GMfmVusPdsKxpcwMoxbZePu2a5Su9oni/Cp3NvdV
5XaZWmrutZgunMTX1s6yL8tfriY4bXNazlOar0dKZ5sUdEER0o0Qy0bwJ35l
0F7M53XeGYYS/DlDivUubNoTR+RTjI9aw5vgSYjdsQoOnLEaQarXD13BxG7k
3l4C76kFKQV3g1/T4KwIGFgYSvu3c6mBEZL3tOkwEBqVxS2NVdfQtQW+JK3d
hlRW7muMzAd36HNZtOOCGWfOpCa0nIIq3lWsJPXbEZI3h9pYiedVfDH9rwdu
+cSOXNZYt/G0xegz+aQYjEmUslxmAVCt9stjoUmry/+Ij0oP6Fvwqb+H1wxp
o+nvrwQzCj7MkBEp74x9VLPIr6BOgGHyEGXmN4I0zO2MP+gx/Lj7CLhg5KHO
AyRBCWmlPbmu3v5cZHm2g/eHyR488KAK5RGUKQAJsyfnj5+/bbuh1DvCXGPc
HmyIlaYkmfd15HaQXZFxKHNkiP9tx7/D26dQUt+OAbmEkFuU0r9tFeSip0o0
XkdXEbQ3En1L2UswF2fW6E2SWpBegIsQ3+KuZtmPTMBYN59TtNf5zA3g7tKQ
NaCex4x8lT2DMvHVWyv2ZjPo5l+jqqy462mzb4bfv2rbjtwQvT0/HdOdyvud
uNdRtDgfYq/OABzPeOjvT5NZavEU87nRXpbwqZLgBcokXMxo0OvBQGAiQlym
rFbW/wPlF9qnY4vnDh2KeppeHyy2p/ewuNf39gT99WvzNGciy4K6c5fJ3p3V
9qouM4BD/3wPTZiufSdFiuLjZmOL9FgVyjUzKBgyT+tZzCnQrgWbM/tpypgH
1BZZPFgn2GhEo8KpqLqLJ/NjUc0zyNGLIaZJyC9RXNiCiPHSALfBZydoUCHQ
+VUMbGbCePRubIO+S9QD0Q7pMJ0g/pbIBoK1wCH1EXWPIi99uPuZPVDBRU5s
1GwLb0gMCejb8EE16cPOs0gET+lK48ctn8RozUU+/cIvssyAAOpXOwitQx7G
aBc12ZzkcUGr70nLHyy1FQUriTddhyWSoyw36IDY0SEXcAeFZZhUYh08eOIq
Bihc/IcfFaZDoJs2l0/SDg6lfyjVyko2tyBBb/IcmaVF5zxPUNc2EYn84dx+
PoCctmBSJrEXVN1P+RhT0JfNptHGu/Xhfjmx7kbrP/9ncEv3BGTfxQds1aHh
nur/S+A7CZom8jXCBy6/yKv+0hKGca9Z94lJSdCFvVIe2bSyDS1+3QyoM8At
jls2NaNDjmuR1Wns+iLz10i9LIcNUwlvPFJwjiYx8fysohm/G1Z1sPsJcG22
YzewNJwmNrZxrnGJSBM5tX6S3lg11f+3lc3d0F5CvNmQf7j/D/L26mIuKx1T
qEgpcjCw/6ylW+RsSWog9rCapAelWnaKW+Fpq/8tuTGI8tPpEMImlxtkZE3d
uD8BOrJ/8SRlz1F55w2Ngnung0K6ibrtFUfWKqBYx35tYcDLhp3DIMHDkWNM
2h5lR/kAiNbhaAQMZfoLhTsu1oOQLlUAgvJ0LdJ7Htn8GggQ+nFi+KDR6keE
C2rH/O5lB7M/lpxyzv3TJGuGWr3PuiIMYBZHq+bwfWPTqWYRCsmSRnEE+pXY
6Ld6V1gcZuEczUBK4EidWtWFkMdQ7X5rvxD2kGuFw83vVISODmU1/Hg4EvCU
RvVvziTuOb8BWrlG22rq+dJsF1pQWeP6xE1+UGW7/29zhRRyZRo7NN9Oo4F9
O+yCrUE0M2KqtrpV8hWeuBlK98Qz1il+xikSDXs+VFQpV/iKFhzTviRlw9G3
svSLhgz3NfaxEgdLHamJ6xAqWtZ0ZbhsPkbbNcwp4qFJ+wNHpSW5Fy1ONC3b
1HbdDIGnM68F6GcpeqVnycirhwdT1edvUKkU0UMl2z/1woLFmQGzQpAjLtJQ
P7eBUM6VgsZ99+7xT0ceMa31bvBVVe69OtgyVLtp219KMIBtfDBcPXG5HuwM
+w/ZyB8+9Mm8daj8d1Y+Jw0OSmWjpBUHqyjxdcMMARTjYOLe4s0q4cy6MOtO
NuQAOeCVXE5xQSB56uWECjBpVo83grtyiHytsCN7KMp/VJXass4BVzQJwTlA
PFv8FH4fHAIQPRBbL7U+2ljYkNx1fKMO0pkTFDxmeCCrD3sBSDUTabHqR4oz
7VLOO29UoFOpZ9yc6DJWwsvnTD0zCHRw9keg9fc2Voa/NhIJWKLhxfDY3O9O
AgTK7oTLeP5NaWr0UcDk+l1iTKN9748n5bm5IFdentnGGQ7X0O2DAdiqjzW/
Y2yGZEQr+MHNBEsXM2uNzG8CJuNrId3JzMnXN/4r7MIkvPK2E7CmlbIk9JGr
A5c8XcjpulSem6TqBkIL9/dISbfg87P3GfL3RDJMpP2dN8aZDVbVGFCiaJQ8
1HtJMwiPoFEExj9YhjZkL1pQkj4SYqzMs1Xhc0RGNfUQgMrj350nloeziGBJ
zFrlMdXgpyjuI17b1Fi/UAq3cdzGJDdKcTFEJjR8hNtp7Ij/mngfOnzFg/6h
F4QD+fAaEAf7FYMNlKD+4xJXU6snDynurwtK78+0TuV1Kyn3lZZY+9TxYooO
EdVlk6hKiWQvMqxaYq59bbOf6EdhpWxhN0RSKVt8fMnVIaqKdxg+ftuOY+v5
Wr8+0ljhG+wOL8S6TDpGwJCL8W4M2Q0WzLWxrf3GjRps0AFqpAO0ho4Z/2+4
nflURGMMWrlss9OS63sKdzuR1bg8wrZBVzZxb3/bfrGToKyQPZK85FXQMc/N
NtlazdI7cwg32h7G1gJQcuI2MbwAcyZwxST238+g7yUuvBOBEdpgHrn9fhfg
0UwkofhLEOeO8OKbdPPmyMqjKnqj3HCbdnmoBto33AdCpIgsqXSq9XsSv0Up
hl7f7INWGQc7dtsy3hwP97Q0WTjDFuhRZIGdw1GoR0/reah9hym960c/M6lv
dr+Sxd0se45UaRn8QnqS3VOEGSWnULI62mWPfklc8QN69UIfYCNv8yDxVIUT
UQ75Nfcrs8cXdHPlI4nyW8aVXq1CTQDKjHF8pCt7vib78A2krJLgpV0R78br
Y1RRyaKdsrtT7LUZBG849AL+Q4TbI7zKwbW+Td+/73yUgc4HUdE+QT0r3tyR
y1xDp+u3D4D5nJzA/5N7R0RVEgz5jLkzGt9KLL4FOs6Sml3y2QDnuQxzQKod
1twg224IeYpYXn9rLsJYztn4zy1hoTJ71J4kV6dbWiP2dgmReDvhIG5+KGmo
KAPBnXU0ICsSh4d5S36HNoeoFdaPQdB5q+IwMol7IJbCh/NKoML7OnYH+La9
cO0BieKwOvq81cFEMmxGqv9UQ4SsKmbllalC5+FnaIfLSO3WxNxGnrKWBHGO
uhNx7OUFuSM52mmJFqNv7NrZWLLQwjmJgbd0bQw0qhP55HReDXTrZEkOQ6D2
Llmg9uZH7iZJFEgkislxuXPEulh+6SEwCK8ZDvHKcsAIaFp2uT1K+5wVUk8n
yMQngtIvJ9ZqT4mdCixLgK2+jLX3zQ/nRlCX0jyE84Y7rC9sqpC9eCblyno+
Zy9qjqA0f6OwiVk8s46OPY/l1t1jqAPu+pMEHsi7/HGJoZmD559zaZ+ehPR4
S0ftyz2Tcl7YwZNkF7uCPnDGXWQiPITvhupclmYb8TtbgB2F8r+KaPWE6vMQ
WPqgPPxhNP+6apQ4uuz6GGmun0/fhf0wOHNUnt56PbtJdDUzOJt++5wKf1M6
Kla5Bu3nF5JL59JureuxvUAibNEKSRRnB8R5X0nXVwcmldvYj1hasbdztrQU
UkWKqp3sVSEeKelynLvMI7wX6xs3J+DwUx74Er4dONaN/jxURii1fiJMsS2Y
obE2nTTZ8uxB948fuFKXKJgeftJW9/k7Pb7eIJ9J78boeaWD2laL+0zuvL3s
CIxMINkLAQbV916BI7gi4wdxXgwIipnluhr8U5r0eLK1kkl0FGCHYypjEJH7
PmbWFu+4jp1tcgVhiGZMeIvXD6w2hGbFAKKkmB89Sj+7EVYqrnGnZPjmg33j
Mmj915GvulOfTUoU+ORCK9zEVptZXYtSAGSrKEdVFL2gsLuue0vxiq3J4BAK
reD+WXlPg1WOI1s9+Prmao4Z/Zl7NoOz9kbHvhddVvXHo2xc7IkmDozGeWE7
W0ZfhRMg3ZnMjI704G4yMuH3aF1E7/8s+1nEGytDm1UJen3H9i6MM1Z3nbQn
EGi/IMHKRu/R6LqN+S3Vyau9Iq1H8sedv+IiX6oES9piegCNdyxH+mcEtmU0
S3mUUrTGp0iBlpEQHH2F1MxaUieVMBNiiYK5cFlcMD/y0l4esq8QUijFnBUy
jhENY0DjFLpanE2V7uQWvQ4mwXAnuJJI1NR4Zm9ey2is1hcF5I90pbl8kyej
RaE7OSHB5x4+vxtVtfFp7qfMh3Ajv2RfV5pXK7myszAmSC9VPAUnUkupdDgh
Cu8vFZ3SCqvMTgw2+faUBPypEg2uTyUdnayOJ4qDz8MlQqOK2MKKjc2SDi0/
WH+GJ2x3kFECZ62s9skNhvsUSQBZHhFGaMbtZholq/DyXtXUYKwn2kuF8jFd
wI/yH66PQL5ROPaH4LmCWg7blT+X+Ub/kSP/o7IVnparsXeKvJxxRsCIl/8R
g5x9sj5yPcwKDY2MtTmRnZ/lQ1DSimRUqdeYcdgPDgZY0XbYx41ybcfDGX1T
AOf17XGcZ4xii+aQ/BCn84hA+RTY02Fz6S7MZCThbVlvL7zzCPZO3qwhImsr
gV1q4B0sy3rOMB0lAxMLFZMRRhMBYxLIg1IYD0JIqBEnHP/YyMUCqpRdTBT9
4mAQslcnoIfF5sgPoWQR7OeX/IFd4K7tGfWQ7oLw+iajppgtpZRLsbUHQZWT
K+ynOMehcOInC7R3v6pyhjPGHV6rZsEjF0alFgoT1QkKNhFAAbPnLzxh5rnu
JPlL+OcAhuca1QMvAw7XHbRmA0WOF31E1FB2WER/RqSbF7Q0PshGeL1eMhBk
+WXjJh3oc5Qw2mR81glRYO60pMx0c3y9wnvsEekdvT4JtXmarQoZy8tjhgn0
HsucPG4kkksAE2lgRHp1WFgThD5vx5WL97z9kZClMpPqaP1j5xmnNP+XkSuq
THmPER3yibxSSNn1+6c2PTIPj0ee42qv+5YHrhXJTVU6IpfgmR38TegVwFC7
Ga7hDL4P9jK+XKF6eh/0ROmR8WHee3U8638nX9L5y8rWDX6dukRzd3H1FH1G
poyywA+fOddG7k445ALZf8w/wuJCijiQNG8FKBUUnB0RwsQPW6dmzMmK4Qal
u+yMqk9q2IJCEGrbQpAudcplgjQ2No7yd+tHsjz/ZCmo7VsnKrn+KYa8povZ
ixOeIvpuhK0wwjK7BMUS8uT/JxNQ3zpjozY3NOJsLrjrCORmM+JSMSjdKYxc
LVYdAR1OEspbbD6O3pXdXk1inBupCEgf2JfXSIuV/fEwXbGGMg3NFPKiYqQv
BI+kiTRGHH6pifkp8BtmwLPfq6TavzLRio0FK5/EdkxKRGWDUpFx09ytUwZA
Sf+s1mE31nJmdFFrpONoyvGONfdMIpYy4+Dw9kraYtfgyvvavHZ9Jv8CObFD
Om7GOLKHW5O7b+T4EuZGwhCAkDihZiWMT2cYM44k79h8M7FWhUnX6LEly8hA
YeT4ecbciIsqRMsyuhRzIqCAjUPmq2foL5r2xCdlVXqc8zOSC1QegYLKvFio
7Byv5NAfeHDEprmUXNy+qksaVb2xMKi+aLHUkFzYoLKtM8DvQ/rLa8Sth1Un
AcRNDGJCOo0QYBx0X0iMr9uM0Z5QK+AX7SlR1I2wkpyumd2rKBnw89NBI0wC
498fI1HQBAcMX3+O3zF76YA5MufJ0nj3K7pkUaplWAOTR9GqkkK1AWuN4giZ
MyONTFJVNjJPyGLRMRCKxicEOkAVL3T6vt7JPqLuPK8jkwYb6DcUQiFzH1VM
i4rTJ/VhEEF4NzUFFGMlvWsvsOFem0x3WdQrOqg+ECJI7tJVtP4kNXgRlneD
mFSWIONs83ij7yWzK5xYc8U5uutKX5yvr2EeSORRdG4wizk4MQHT4tMaqQkB
g9rNtj49ZxWSynns25ysNBion2k+rr1glGeJI3JsCuFLEgq3qgADgiNXB975
oWF5QFKsApmilcKmwbDi8tWYpzKuqzC93tq3W8J9I2hu7spK/46NYDgVAdlD
MPyLHjKidskInu9a71VSWduJfvP4SesGsfOGeSi19bDTVL2GzVX6wwvLKEFZ
MYa6BrCeFWLPM0HHDlqGbCoKHLGs8NCWO/iu2M/6hgheLdccN4wG0ZQV81Z4
Ep6nRhbVY1xoqJsxuE/Ny1tBb2f4pStBMpQu/N4qy48DGCI1KcYAtUbAoV10
6lbTiTqkxYWxkSAAE2fwRPHnTORGCzb3c1WXZeDSWUosxqVGFpKg2W9qOdse
Lr/6Al0Lmt2w0gf1X6MskutukSOznw9IGBCJm06SoJo2kZ3cJCCc+bY9tvSg
owATn8hXMygYk6VF60kXuUsEjm7GdTnuGk3qcRjhXQKQ6qsu+3stOwyX3iAb
m4/tsbyTDQoz47eqHtrqPe9Yd5L3Lg4D9FGC+a1ERGY0jMCpMG3wGb6p/BNc
PLoNPKHHGZ9y0Di33PVz2fUnJg+lEsVlbGcDDQyCmLXixu6DVhgHqN53mHG/
xH5FnLF6bVWXIpacXK0GkjHUetka3I7ZTyCefccATXrb8DL1oiMVUWjI2E8Y
XGpwcMnTItvR3M9r4HRXH7m/tzba0JmoT2Y7PBrYTb20t5MyXt81uegll4g8
WSmU/JRKugblokmJZzkKZ4cIJnwC3EhIdz7u2+5eXnRWTTl+vjzJ4fXE5O/U
rwH+xfsdGz0EB+m0rWym8RCYhMvEGRD+jOtF4yeMPP3Xv7dkEZTSPaZhpjqT
sLifSq7NSf6SdqQcEHowOb4JoGu1ut1V/tMZ8jLyMY4MmA1FAiUcJNk1E1V/
zLWsOz6NLOIrIBbrscx4biidnXS1FFiZbn9Iyoohf29OC+PM7Q5mazqZBe6N
jcHn/07vg+oPzmX8UxVk4irfYveAqt8sIdrLUKIPeP6cifmyw5u27M+VpP8j
jLCEWPxPyI9ADr32gSl1+LYgLm3NKdXa1lpaZt7Iu7ry4kb4bgNQ3o9o0T8M
REfRR9Utnj/SUgtSj7RYVS9eyYnqd2utUio/XsEh8uh1m7IvEL2B1tNSsUIE
heBnPWmcig8hxWfA79qV35f4NpgoCs3IIVFH/7n6zIt5vPQo7dF2qMiIl3kL
eYgUm86Xeergbk0FK/jRcRxm/G6b4/UX0Av5CpHZZIKANZ6/fQhFzhRUB0fu
jDM+iRHpzC7VG8Ore9dCI80Zb+LGTzioifFhl62xFLyA+Ws+G0lqYLn+v4oz
dJRBHZnESvBk+gD4Og/81VJIOfyqDZa+1bnsOO+SWIZzoRopHBSYRlJwSFS6
7jxRkrW8ZpoL0SYHPP0gpHK29vRsk6Qf/b6BMkq8/ThZBMloJnLsuQghlnFu
D1/el+V2AVRUbq7pmTGd7KA9zFjBvT2bU1Sk/L4s1d4x5jh+z8SljNmAs/Lm
6h0yHQBrE09BvKbKpmpRkMGtNU5Sb4ouaQHybBwOhEu7NyXxPhOwRGJYEowO
B9/ycyKHBB5PUSNU5th7dAu0Zx/BZLFU3/v4yvQTOFJh+XF3DuX52NXgnKX7
ykaUoWwIHo4v+0tounYnZiMgcpsD6XBwYpQUCg8DzKjjKAGIRHEsBTXCDWPO
/eiVb9Ems0lG1BlDbLTavJIxJpk3j+a1wZo8h4QZMNnqZgxUbaBtmg+E8qKU
BHnmw8/ZhfDs9vCdzUNZfEZ6OPGfuKg0zmRqtFULDyuE0A/1kJ3EKFDyPwEn
ASwVQs7UlIGnLOGKVGvHF4mNjGs5r6K77lG3P4diOG9VyI6HjWYHCmIdf2BJ
CPBNzFKVOVfmsyDpgPpb6bVvJNz1P8NCy+gMEU5Vb22a89GNGcVlio7990kq
LBAX/Myxp266GzViTdckfVTlqW4ghp0ZUBbIm+ITEfguTjkSKNVhWGKGyvPE
Ftr8yQpsDXiZWcwl5Ws9iHchY+QZLzmrAOX8FH+iBr44tpFjt1LZ8eiUL+tY
BQADBCzsfeg+y6axwRXQH/plVvQIZlUepteJDFhQjOl/a/mHN7Wam6mfM/K3
sM1d0fuGxBxaSE3BVmdOpErrK5AHY6IpEYbQklRoCRNPeqUcj4A8aPky1Piw
0R0Q4o2xKuIo2NxAK+UeuqxBcWAk55ptgXG8I2bZrXjlubXdogG3PZgpjWJr
QdxefAvzTiCbEx3EbrsE0OwBjvxPqzGx7+4z+VHtZONWYgxbLrVVTyaSguF/
g1WzrbS5EWQycokRD4ae0uOyXIjU8STiQED8miWYr2xmLDPOlokUlIs9RNgZ
Yse/B0sjjSOeNH7stR/8eaMogzx4+t3PSKq3X680Tm+OkSTFMSGu0ok1Tdkv
sW3DQLoGjfABaBjeA7Bs9Z9ZNCKBnwDhqgLjYcFJmb1mi917Ku8PaKwxAyRh
Z8Jhc+yEb/MwNUtOSrVHpUnQ5YbHhEi9fmTdFVJUzybB4o8OxXJjTRoTDZu8
PP8izwROLD4EqjwrVWJaXbgJfQs7QDgo2WlgFR/DHFUmMJazd0WEVx6kMx9G
3h2GA2xT4k1zS+Avvaa9sPHWIDwVICvIp7h/MgqFIeCbC+za2m2I13F7ImQm
py7d2zeXgCd5irwfQdmEmsJ2+MrJr8XiVXGXafPv4mjmnY3QOdEhVzAPyC8u
2huujfT9BG+SUOc0wnF8n9tybYWWNf2iOOLfUUe8qeWlJ2KqH71jhniJnZ2/
cwSCa6tDysQ15AV306tmlyXZ+U2LpYbfC7tb7aLSCn8UEw9Ztw1Xx8qE1Fve
Ou6z1IuY4zl4uIXz896rsdaXGKemJG2q1zfqfPkrrLOXkSC3QrlghhJvFd3W
37aO5zWA2txyf8PdwdoxKvi0miQ5o0LckPa+rc1E9dYqcrwXI10HRKIKzlnK
DvnzMh2EFykbRPFe9Vvfs+ybX3hzyvF35Qt7/vu5zE3XQCzhFwpoz/ba41yf
rLt6iX+eko5w1Sz88B0sZytLI7f1YnnJ/sFBfbqftSquvbUplhEb6gw6qqVt
Fcjnk5+5fKvTukzNcMUng+84DlzrC3fDz6+C88XcMWHxDrSL+C18EzyL+6yN
LpJY//c2QPlOEBJFQXCA3UatHM4s9jhU4vggYF7PeQFG+2beTPkuqxo4eJ5F
7UCeiuqb0Dy0GKeTORKtOT0gYQ8vSMlQz/77wuPf6PLSuIfNmDY8yoCXnOpV
V22o8zoQDCQb4VEnKHSGj2IQVDoSoK4YE+3vg/Ni87fnYDsfLDLJjieprepV
+cqHchbU2aKiEO61YvjNYNIkeYdcYgYz0XzW+FWwLoh6Iu2EMrsJyW8Eq9h/
wO7Tq1lG8dwZeOJLo3n8KQD1KopufUxv+8UCA/GloIvGfhPxnwxIQXijpaD4
SBo87oyGyfpTOb/gsY6OptnvpoMCwVCX6lE5Q+LAaZrSF3qbjzI5eSuFVFIH
r5k6SmTokcUkzw5QsKqo7oy+Qi65FkVtFgSSbymN7eaPDY2Ecrn4MIY7A8tl
fd5Uc8GJ0+f5VJBuS9bLpRdMu9biu0a4oaeqX6Jk46yPA/VHVrY7GKlzEOly
M0MdOM6e0aVwv0WDDtsBUIatkpt0e6h96RWjE2r3WmCE89KJq39xm2Nrc+Ye
nhZY27hVlFwmw3FeAT9ofVfR2qxfpdcPE/egy3vHUvlFRjcpQ2S+aZ7z3K3v
nz/b5if5ul9rgcMe9ouq2ARl+rrM16/nurOpOC3Af+CdIpPDB3ORazYnYG5i
ygsHlr0fAmKxRzCQR3FUz71YH/GfIyfHv+Z8rtNWttDUJDzND23UmGKzicNQ
+8nxh+fheRYv5Cn6DheWILKDgTU9n6/VS/mp+WQEoydqwMhaJhPLqCZAF2Td
Ldit9Fhdao4wi5TxeQA3lS442fFIoAQDd1pNpm7pZ7qGTkbmDiCWevqLlbR3
Uy1DosyaWNpw2cAieg0ggEY5Q1vgiFWlIXKH37g4mvOznqVrT+P9t7T68GWW
JJtj+stHpG12JYOKfjFd3mXny5nGxk3dI+sqa2pXdq26c/IWNp5aYY4Ob1Xa
lC+5kaMa6LqYn15aqSaTAVUYLnYHzmn+m9Y/rweOlWAqydSW+tMFvI9Tvxke
9Qx3ncqOYBdkoq1YW1aLmLjtIOkZ50mO9FwlZhkcc8pIbwuNQtmJTOT0gZaM
wv5hr0k6IxZq7E7DqybHKcbrevDRB9XkRs9aVwb57buCF7eJU+Tb3LEXHw/T
hm77Xj0I7Grfw6RsoqG2m3p2nS451GRXAGZM31gxcDrvFGFTE34YtrY88DHZ
Rj2oAd56vQ7aWEq62SWebjHphyCRpCJpOtEZDEt4m0OcgYcqKnIwEnZNEPk0
rMBqmj+6glPiSzEfTiMU+WQQeHPbAuVafYO/D12a5iYgKhJJqfIgewW2JlZ2
02jcTqyKHGdoDP9M52sTaKiMbZl40l1OxrLA5rJ7enlINpumqXoZyAJqidn+
l/IzfE0GsLcNt3EOSMd5nx5OB/1HcjZlGXwGufARNSQh+mbtlPmY7nxZG0z7
nju2KUEFHUeICEfKJuppJ204vWxLOh+W3tzxlU+6INIa59R2HG41diOO5THM
Ke8lG/+jJgRKoBrT4Ypeu/lbJGaa0VHq3QMwDJWBt/skl0OwGF236hUZGHpA
RlhjXZJLdoQNatzWiN52+kGwIFWqYybIuAuSw4Jn19M8MJztuSSF6dWrk40o
PcEFe5UDhRK81MvFQHg8WY5mE+OLKSFE/Zz+6Jlj+gy7WAgbeynHPLN91WLm
4SxB+cSI7ayUJb9fyWxnH3bs/2OueFgoNKMPFEUDIY5BeasYHyp2k44lyqnu
qQ86MYEvol1PCrX6/cLq4gMgDmy7WXwv3zw4rLOY78pRRLxsA0H/XsAFDvDQ
Y2Wh/GjXo0HcmAriUrxPt46tsDvVdVst4dMx/ghuIZvr/GdEznk1bSA3G8s1
TGd2FHaNzAJbmgyHhLc4Id38XNegYTT+pasqlBwNoYmUdGywtKdKF675mLJG
vnCaDzlwVWrbdrTbMe/XQFo+i76lNBa//UG/zwzA366y8rhr3fZ8IjUZ7h3z
iU0Y4KyyPF+FFSzPbaU5ssI73qSh2gkkgr/496Ww8IRh8KbtfnkILGlRrWOY
9/eGBNlecKLyPn25ykmelUjiZ2wlGDq4HrMHxRTZiywz2/wd6yxpDNy3tHI1
zcT/2ybsQiDTaBNTkFGXGeMniIwlnSkMFuCxl01TAs0KouMMxm9TLfHLfUuG
Dwsc6n1MWSWzhphXEI8GV+JYoDaEqiuaGzigwTiKzo/eOQuIf75+qrd2BEyg
Q/Kr0ykfRfKUN3jUCNeFV5MWRfdYoCkGh3el3zmcpiYdC6a5VZ37q5XrA884
SE2WmDJmVXrD2Sh5TA4k0iIK/LjqbGDZjekB7STwtH/NtVykihrW9j4/NNoF
pZ9by8ZXdG8kne54FTsLmdoc0g1RxmFfRrQ2tnocxFj6kl5OZgMOg6V4fAIw
vlpXw+Zm9MJvr9vCYVHXnE+6VIUPj/cPH7JGYxH19kriDIrE9P25O4s29Cba
m1nu9U+4Z0buWcxA2J0EkKTl3ppk0b4cObaI8/mvK1Y1Jb8/9tOy/QHMuW5q
YvwtMLl8SpkFffD5uSfRZOfA3NmSFp0MNoZQhYqcoTsr/1CleiWViZfEYBBt
K1FQI/vy2i5Fs+EzHqIec2ogIePhCT/1JCA8IvxI9WQ0+NJ0L6qYo5kf9JZ6
N55mHb1YfdL1/B6YBtjxe9S/9Eubss7O+FKcbPwpQdpTuMKE3LnzkzKlVvpY
WVVGNpkGTvTjVbDDWsqwYke/ium+O0+gv451B8GmzL7JVoQeyXs5baFU310v
p6xvw6FA/+ac2Wf/8XxOhvdGJ7WYcbaSUv6Oectv0sPTGOcWsleDb7TLooKg
nc140Su5mw2976UL0KYoLmx+0FGcrJ8htVEiVg36Ubq4A/4rMc0NzuRIBr4Z
dsxzGTzdpoMLjx63YHGFxHEi/KBKbssksM8BqWENyHQtLUKZZ13hNfHuViTB
VV8Cnv8izPwA0w+P5UQsX08Fn92k7NIm3cHrIpiJawJMBMiKJQ6/BvsNB28U
Ci8gcllC3J8hdfDam8Yl7lFyucUOG5E1xPTgmJkxEEFWftUKijC94GrshzLT
iMp2jN2UH9uQsZxiGv+ScRiIVdmbXjeQ1HVstB1WtxHUKI7Q9iIQMplJ5QWV
Pez/D9bIFCc/KtEraSm1DuJyp3+NwFAoajjPMY2fptHFoNwKRJ+oZKqKbSSs
Y9NdMu+jB7EaBvDf+Dwp+XDPaNUkiFCiWnLhCS6CfZCiHLX1G8QkUdKUL89f
A28Jt7xn8N/zS5eHZl2yQz6Y7O/uRubkm3v4hcmxFyd00CC1CrxcFQUDj/4w
3JSk6PxZzVwWK67mgFX5MwV/46p9SUv+yPhGtmEO2hgBAf6dONXpjYuMQyYP
FzwpbSbKXvLfXF54g1saZEOy3a+rhXkGtVnaexweQz5X6TiM14kCecRJFkYv
g+pavGfvKV1kT+0tq9MXdP6oQuc3ZNsu1bT8h4WlT5rc2H6ZSTvO40MvDSGE
w4F+dV1C77fMJk/PYQ4JvrrkGeOnrrQ/MTWd3qWvXtWHLdRa3L+pqHryZNw/
QwdGYDK7Nz8Ut0yHXFSMzcMqkSwCxx7kx+vNVUXH/wFIoMGThqs+4dhSTDU3
qOQUdJzBelM4Yqu76OZ6KXww68hnCTj7wedNAhGZZTY5jxQtqT2gk8bqzvuA
tlJCR6Z9mi4OqrKzUM1DfBnfDi+l0DMf3n2w/rNnlkwM3ZZ9XTehJDJPfXK2
d2UUX0A9kPwnAW366H1RN5HMCYUIhdtTiKy+6bY41BDYbut2x/Amn9cr7JTS
aTdgzNVd0dUsB/e8wHPBHcwF0EmmoCwtAjl+36WX8rP9n9O6hrI/XaajWj2Y
Fj+3/QklzW78zeDwKG1R591BkD/h3VyAsZfVTNR2qg3EN0VXhw2CF97E0h8Q
zCcvZvveF3xSwGOD2uTH7bTuN+XYtHH8fBv4rxg1T6pnkI3up/DT+oFCYysX
dWv6lla45EP3UBJsUvEr5IVQL0UH4PNuvEtUbJjGhHy8BJKKuuzoiCGXwoZc
/PLe5LKv93V5NLUIyikrxgdT/W/b1y/+WMuq8Cp8EKmkVNs+OFTPHAnWCEXz
C+2qUsFquqJVe42n5y8WHA6F6jblW59JqMS8sqUcWLi2pSNc43H5z90wf3fM
EeiGFXYNimcOq5MT0hHSfqWGeSHnNmnIn5Ul520eAuGYEAINUmCMFuAdw8hC
suBGzeT3Ki9LuFkIHYyHGb4wbnXrKg5oozdva5H35/I1ECFIRHVcQcUWFyMN
fsD6boiOLb+nlGK+SNHJeXcePeFK4oMKOPCxp2Ay8QSiSL9SK4wPmM8axF2X
KMoqbVVoWLGgzW8SmZH+XmI7GgYA38XD6ziHl37AJrsnsZ6skVqXsaFda/E3
YCW0G1ht7/23799tTQKiX8t+M50RIvz21iVr+gPWYB26hsJ8V4qF7ctZ1fYn
qDE8ONPH2TSPe9PDqKdSB/SisDszyWdr7IxrAscTMakwzpPhkj2j7dNUTxvD
dwxYUmnqql8sTs2tle2r1s9natg4wwxgT98uPk9WeXKEQGXvhi3SSz93hJ+i
tsPYJzaxZKvFZP6IZZJXU5uM1JvbSPbUXSRVQ713RkPnh4x9daLQhufT4Wa5
6SpHihtSzZcmp2KJFOb7PrlrNBPnNgMs6bN5+nywu+ChPKzSvOcHpk0wa8VU
afZJEguI7EiYVoa+O5c8vct1r7WSr/1EwqNJJ0Iy14G0iKe35d4Oz4dJowA7
09Yyv8eeADPtfpnnvewKuaItTs1oxgFl11KFY6sQ2SqvrecGZVk5xdqBbtxm
lRkcTEPHH+fujr8Cyoaq8zTGmCfZ2TyJt+hk5sutRD3aiWqLDivhlpEHg7oV
KNhbe9cv7TrYwy1Ln4pkIVWxIarbDRVxzoISDgz/9ghzl28EPosqtxr3HUUg
BDao61eJWcjp0pVu+MU4x3kDcxwjPMw7hJ4A1t4idf+vemCRHrjbawVXl02X
KEYtCO3fEcL2WNvrZWOmZAaFhM9RuhQyk55emQtcVOo7g/MOaGQupe1GGoFP
QB3EB+bKNptRK4DmDb1n+zh6WCm1g/HfJw2cjPhwfXoDiVrMMT9er68SE/ZR
pzvm9TFgBYIFbj6vzmb0vKChj1lRHE+setqAchjSxfZd18d4YabULLbprnSQ
z994JQL9HyWRKbMbZfeTXRbaqX/vVW56wEY9b3VmkQ4wZK5Pag2mvYKM9lc/
5yEk1a9hj2nqwIAkSglm3YsxzE9LA4GZXob73BujyMtg40QJNvYN/UWaQng0
+9GhofpkGHhDH3RfbnggPFXwiQECCQ+Ed/Yi6nGiWGHs+/JcuMIWI3QCxKSw
qXyGVCDpGq+BdRE/na+aQjS0sRbMHGrtm6u+gYmbd1BdZNyiNw0ivOr5VNqi
boH/mwJBRgw13B1z1DOWgv4vWw+B4HXitCE+3gue4FvQroN5rs6FtrJ14kgT
IrIRztW6//wsP4v8tnJk9X780hqE6GroYZt7N4K7chk9r+d6KdYPEWoFzv5k
Rl+/qYcJ3WtRAincZetdApJwSQmI3eo5yV3lSRDcW4xGrEJNEfEa7ZcqLuLi
R+VfFJvyhig5JajAqZC8tqnzizwxz0DqRw8o779x3XdiawfkmLjvPBSd6Jeq
4TIhOks8Y63p/E9KlKQzRldWDRSdSSKhzFh+992h87mjpYXdBJmHw2Btmwl3
DNtNW00Mi5QFjIffg4+TAzgIJDl11/6pukDmTl/VIBKzBEqIy9q7lGGiR25b
rszy/CSRLkc7SgyXc3SicY1pSOf5CsvDA/n24TqUZMtRGvyyyPTPAboGaopn
iXeZ3W+IfmcOKFCLsefoNS6zzWND5oW3/mqmnc+I+7wpT4WoFeYMajfN7Hkl
vqbbGqUbd+aWZB6+Po1JoQAa+D3fO9kjnU2v5hdh3RaBeavxCwbx6ZowiJDc
C+eBVRk8f1ozeWAHlTBalqbpCHM1+zR3aug/CSx8Rk2sAk1ti0pRxbd/Meal
M4DHTd7wt3/ZlhMZUJ9V/zknW3h5KiYuh3BbuIVcPiJKBx4ReqTmV7hq30WJ
MRTesnJdVv8Nm1Y5x4ZNVPXrnwjtqVsFXdDRi9lipbvcYUp+ct05MXiKynWv
yQ0FS6Jflf6d0IyTPsd5M9DEZESz6ZrV/ZJnpA0GnvPa/3K0JZ1jLhUdvqo/
XM2tAoGvqcQ+I8E3nMg720dyHGpJrFtx1UvyqfsU1rE8bJSqNdD7ZMaJv8En
ka2QIKXDTdB+0TXFt3ALbWx6wK7xFAQRuoM0QLh6dQ+fh1vFPMe+mPwtR+uX
Oh8vCv146TYYVmQHWDbk3rxXiOXqL0uDuNalARklMvTxk9lHYoc0EXFfFldl
3LjFwva8jx92jr0s4PlaMVMEyc7acg6uZ1yyQ8ZUaU5/ZrhiCDLpQuGe7yh0
lHkn6b+zZTd1iJYafMF3OcTtz863xrEapIa8SWFiwlf2LA1k0zzbTdR4eZlu
9aoSekL96K+Wv7XoZMDj9aYSR49Fjfeh1+RI1mDVeQTogFT4+jnR8wKtygxz
Op1Cx5pQSycDCxcUGOEyKPgkjfPqNWUgr9+RJNhetylfXn3rKl+pZQgMk/Z2
cCehLsRX/1kwN+crywXKcxVU/kxwnhDU/gZ3IiJh1KTUk9wwW9ty5FBxiJl3
dDZZbWpLQKOF5kKBD56nt5E7sOOFkXX9HLsQYyaMMxevDfNcnLairr3tuPZL
uXOFwh9PDB6gRKah4zAdL98srtWb+1W84EPFTeM8DkIbpzy5KMGkAK0udto9
vPv5bO4wStosr7xavfId1w41yVPCDSS8z6J5kUJTmvzStG8pYiN3uiIZTSc/
kaa4CA/Yq9juSCL9Eab6kJoDhMRfTyzWl0ABpqm5d1lAl8vSfjYhRgeDHDeH
m3P2z5W6QpQKmEFVQoPiNkPvcQ5HZlOJ5sBQcBaT2kHNfCnoYDgNwfRb59L4
4hem0QF/iCFY1uYYatOm32j77oD2QdUTjV8qFNit/Ci4/Hdq9Xi3c4Kp8qr1
oE53nTqUCdppZ/m4tGfuHQec+AvNYaxu35r8LtnerqvqGC7B8WQFFrc9uFZx
bCjneom5jHSHiooY+hahOJMkNfAe3Wu7iy+A8cJ2xo6UQmiLF2yQWKVXvz/D
P5CHw6hkTX2OjrOVb9z4OlPMOtgTclPMrJ/B7iW1pbznsxoFlOvVlhGe8zke
Ae2Pd1qLY/4ZWlfnblIqkNcD1BMLl2UIOk3t+67mh9FdolsyPrFQJQNInxI/
0CTZf2bqBtz5f0qE44n5gSCuBWnaI8CQ813yjkWFdj1RkU5DdaoR8DhIUYJG
QreWCTD3PFZZp3PDLk/wCaGmJHVzUMGty7gvXXa+Mtq8SaDrOBj1Kygf31NE
p909Kb6WXEOR3QVkK7Je534VHX82zAdjZB3rVmlbkqSbMuQwJCe/A1v+vB4J
3Acx0qQPBY6a2gXUsusRHEBB65Hpu/SrS2FmF+AhSLoQwvFvznrLt/iixrQf
RssVvOQz/xnnW6o3qHIjvkQSfuzsPiiEAxMclANCpd5FKBNUW58wRTeaKg+E
mI2wzQP27lDubCgL8pvcbYHqswnHUKbnzfXkm9gV6MFw6qfUj0jAmROu1cQj
Er1HNu/7bW7WPQ0ykqP8foG+fytyrDdo4jRZsnT5CjOtGJ2pZ8e1AtGBwPFK
69n6BHIhS8H+sLpdenQuBfke7wIG9xBGgp/u8BgtfkuF1T6CaqjDV5gyw0eg
HprWEAr/J4TBWMoqa8fF5/7tA8p6geg+WR+WyRCb07G2j0/oujIP88vnGMBU
qaqpaf3nfbDhcFZMcVcfODyOwr6C+gdP8SZnfW8KoCPXqhGo7/YsGBRVjkFp
bTyjnw/lycefwgGY0+gTgh8gYdMM3N73jeWMGyKcmOzPBBI8P0y6vzIEPcte
cI63qPXRe2D6uxTc75Ko2imI5DXFsJ01F0FIBXZDsvlq+Zz2s2KvNDpHP2D6
HC8th0CaDFUWXozYx3GMOSNgf5160+W+5vOEIqdY8pW6MphIsPWtlwW5YIZZ
Zl74yvKXH+4iaCrcpS+YV32bJtyS9h6peaJZX3i/ppRwih9+juLAyV6tWJkG
HyCkZnx1Cy1HVODRJGvnVo0wALR0+8b1aKPYKh8y1luYzXL8b857V/bq44HX
6SDpjFeX9Db0gsDHO9CABugdb+ZvAw5DoR1pOpk+YBQ3xzr+lc3jyU9g2P/r
5hkzsVuU/r348G5Kd0oCnOhJ4iX2BAdV5l7KfVzOAXTjzUngBgnWpCZpqksn
DHgBuMV8UQkhnxs8X5nWzdxe8uBbtlcsJ/Z+YeoZ1oN1O7bmyoiiM9yb2jQF
+mOqnI4YnBWfGuxyoUwKDgShoHPb5LzqzmtiDtKViFv4lC1AJx2+CWUtZ/6e
GAOhXUWnRERgmEdOTPPWkSU5exmFt1mQnMZGUeDAEA0xPu7i7WfVgLWnz2ZP
Y/l3bpqjcfwSNWC2v7yy/Gx7MOe6aCWcjU/QCvpsQj6pxWbvGF9frNy2zSck
rGscMkyqEjWrojgosNnWz0h78PX2x+a7VclNxZz5MX3q7Gl+CWfxJkyNUDvr
lsNhotoSw7aHGNcvTl/pQ6T51RPWxT8WY+eDXoyB3t0N5tQZ0v44teUhXs0x
xdOlxDJf/JBVOoFWgnqyfzieA6+/Bt5E6RCUD+nIqLFix6/gLcKYH5ji43h7
JCIyf/qDdLfdkcDCWR0XJGAcP4vv0Q2AUTkPpMl+pu/Calv/oJvfWwjymXrZ
SDeFJE6YplONVnzN5hfi/7wuiQ7c0CeW8f/+9uyhgG2tyzw33AaaylOFJ5JF
1sbq3QyWjHrVUZmO8C9s22HKWZ+/e0zih9T00jQZxD7OoMK4TdrbsF1u5lTW
KORlJA+7MLWFQS87qJhKnk2dp6F453YPFQN9A8XnIAHKu1BHbpLHY4WTxCEX
mF21+lXB5yz2Vry7wXWnnOu2wJhYrebjHGCN8qfrm3m8ebhpcQSgwkJ/GQ9Q
ZbviuLwMS1fvZwwJAd3a5BT2DteKEN9pWZB+kyqQIPBCKmOOT30SIkApjEBz
U0p8SskLZUmvGMeM7D5YcCPdVBhxF5s+YmGdswTPaxN2zVQNQxxb0KqdHmG1
cnCNsmM6rpiuWnJVP9q9h+hdvq0NsAWL8oK7MRkEkb8DLfFSGwX3A0LgO0XI
H673t+pKV86jpR0i/VLB9yMa9iobUrZ8vof12q/MJuhcnO49FzYWFNLBtLt1
V1uiBKdKIrJA99peRN3e7PCMhK2Aiph0Nj0ngrnrnFK6BOh3HV04AwmKxkbc
XsxFQWzfOhumI1s41KPZ4pSo2sfSM67+ozfL2SGdGkS07q0P4Ayv3+2FjssO
bS6S+Oe9gBiL07Hy18oMAl5pqumsK7o41wdQO5r9YbFa0V2uEq1d+Dcq3iTx
ATphZM5omB8OxH1rgqcXvUWgTAFznNvJUh3avF9Be8p0k5zDBaeJxgp/kC6R
2bSNB1MknPKPkJwSAr8TPecfY1z/kKD1fiBPQRBrOlzh76YlIp4KtMSiXX+C
R6y+B4e4/k64xgIAF8DMEkjbuENSOMX+c00W20eY9Zo5nPgz5G8IgVbyCtXe
aV8q1Yt5sk7RHFMvJ7ZpC7DCpSM7E0gPx2qOn8dedueCs3Bi/FRJ1Uvjigfw
ECdgbyE5XUi6nzCHpTRZtqk8od9oYnaRjl3lTDvha2Ish4fXslLrS0qEU9PQ
2jIh1/QxdzAT8X/7wnULUwbtImdlcJMlH8zGzQN4gsJPLTkv70ZumLixkKob
v6rbcGttKvTIdFyfeqFE1ksL8z59g0MdmHapCeXWtwmKmMU9/ryWWSn9YDnY
mTMyKtbmHg/cVJxVtzQy4etYkdiV00zTGbjZWqRognzY+1yveVj3Vk8B73Ku
fx+JiDM4KpAtGEon6Tct1fVgHDd6Hx6odANo5gwvB1NGiQNdfK0RzfVLv4b2
NYiJ+HsgKuvpvl09sgTopaASjCSKqm6j7/QNiRyIm6YIZbaLyCAL/qDvBOhb
jkMOOhn2XDONh5z47NF6bafCh9k+wwb+YPBxD6bn+RNo0g413j1Flf4zgLLp
K62f1tKGHLw92qHftLyZkpMyo1/o3UoPDhVFiZsvhVarejWjDw2/G/DnhRwn
5S/0JSAl+LijqOALD9Jvf6AKiAV6cAXBm2al9yy3puyEoNa3mlYYBOWcdzYW
flOAoOvWpHzOrrtWHR8QDgNyRtQsnvZeZdLzLxKBkIHLZraLXCcgY+GOBO6B
aTaqIAVOU9GvfVF3igezJPzKWhiOSRmnvDvGCSJFWDDayczB1J+trMw3ppg+
vWlIvdtywQ4haMJnVWfwkLI8fsDWicavFvQBQfDuJO/1UlQbHQsT5LcCGruE
2Y5/e3ZuVFfzUIbpHRANNmOWGqeysibpqA8nXZKObWnhfh3qjn1ah/ji5bCy
rR9xippiF4nyp5w9v1XJPgVjDIbvHAGyTeAZxSD+8PdFoaLuEwrPr4yJOp8n
wI25OwfTZvK+oAjWsR8492DwHDr47bojUgKGqLxnNwhYL/6vDKlSmcLlxr2K
BCLyljhbG9+SHRXV08QCq6ViC4RMrvDXfQ5ocD0+MxuvPBlW+8CY/yGu/49Z
o5MvJw9Y8cOEiuYhyDxnTHbRLXzFjtwhcZYwDvVgh3iyf9+yXCEHRuf3dFdw
jsLj3Yl/A9lmTEGpgW/HYxs0Iw+Yoy0iMYDqUZPytkYRor5KRWySX3PYhhfi
pSGSF3sk73HWNm9ImB9DsP86tqiFKJGVPjO682YOLiten21502K3D+9KFENc
VyVx3gAgKGxjLrEIE2LcYglJxfEG7N+pErrjLDimaIMS4Wuymgo+t909HlwD
Nhrx0LCHkw7ipwxmUAFHwSaHBSUIiQfJ9DR7H1n49Yh1mt/Khbez6Z7RSrxV
wY4kYHPf1dxp1+izAOdGhzhIjSZaulGzbUqoXVLuY1F/S1pUUclH2CiT/VC1
PFLLBd30AkgrrX4KoDFV2oBdFSUYvEkbrPd17z1A6C9Ha9SsJ1KVS8yhmqJS
/S5+Dcf9dbfTTn0mPwStqSy7uYaqwPW35vwBK4oaGZXBPmjvHftRCCsb7wDC
r43e1NwolmfVGzc9rFbRhliUGj86PVkYnBBydVoS9p8ch/WAbdP6FCFLQzTy
o+J/mJR95jECgD1XfOG7v31sF7+PsjAXB8i+QsQd7pnTHx/jL4JdyLPjmCo0
0tydjXXrw1v35nG1TnZkStojmW1OSetddiSmGna1FeqVtevksgRr1hU0IMDy
wOHRfHfg1ZjL1NUXSbQzyj4ROANhaJ4MPWwyVsX0WK1gdyyyArz3j75Z4LWd
J7TtCmC1XsiC9c5dwc7giX3kgiS9zt8MI1sOm6PkUpWLgfUdNyRSGlSyPA16
1NX/m70UMy81EtgIP1VOEv422ngx1Dd+QWwYu28tyTaBMeiAoS000LfCrS5T
Dwy11MFYSdWTGyL5l5I8RLhB4pugPh3iipr+YN8GERFMGYEURsGFa6vhnLq+
a2/urUROk0GY2JN1d1XnST019Webxic+PsVIDKlrbYKw230iHNZCPoypm6mc
JKFEEkMg98WGAopIVcdzcEcq5aDWiRd8fDwrWgdXbKf5i14H+BGVQOiqNiPw
95ukuS8t1BoArlgrM7vTv1w/jMB3CSTzQ3sPaeekk3qebsA0/fyMuhMF7IIP
9iYutbyvEk9cD5iM8nZ0O1oNZN1OQGem7ChAc4Js+TK0lGWs5yFMBdylmn1a
8++a4P2CHoNtb4jcl/3fwxUbTF2FmZe82LjvYd9IaFUHjDcnHVg/fSiAmlPz
R4R1QyTRlQLU6o0gndl3jFG5fl4uoJoJeqdiDqGv6o8oQMcpM1qMxrK0IQi+
xfV5LE79BO/xaWidu6jKgnyyuRtPlpZgt3JYGZCCCAYUc5DYcmElvflxNY1n
rZNSKvLj+4cajpuurbcLlMZDX8vsBdI73WpBHagBNqF4ee7/+54MWu+naKtR
BAoZwC3gkCY1dSee3e+zKieoPDuG/OOZCepxN9ojGlXr8fG3VwcHf1DlENNr
iSzHbNR3G7eFp2ojd+plQDn2+neoG5zX6GaZyqTMV7+wA/to6JJIpubtCByf
YFzPUgg5/2eCBm4bv+4IlVpJBllqZysN+e13/6SC0iuwlUWDMTP6oqzZu3XS
amcmuoyRFn7yDGmvcF8ppU/p2v5Rlzyq0msZ1hSXzyOIy+d89orVO/4JHG/f
jhXsDzz+lqBI7v05Wqd8MFsnP3kynxebhNrqJqy6T4/8PqIrJzGscGwCBMZe
WSigSrJMN4QHi5lZR3KvB4QuCdbOAGxc1/XFyCTctVuQmvbV+NqqHAvUXdwh
E0hgObXRfH1td2BlJ3U3N4+9eeMwaDtfKLWw5UsklQyQ8inkVycami850VjA
PCzSZlekVLwEo+Cwq8QhA4xv6NJuFYAAAeV5dDoaz5fyJ2oafg8IOUj8m5OL
yaXCVnIpg/QNcw0ExpfjpILRYRa7CLFiA7elYjW1i3CYpdl8vQImm8ZCyTvq
1FWQ5KYJfBDXm8wOLO4WRJ+DxyjQYCWolgg4rqd+E6mzhPSP1yIvgAw/pdWy
suC/oxawsa8RzJ90IHsT9h44P7oMj4usO/yrv4J480TZ4ApGf9ykVGk9VJ5O
CfA4Sa7YKC0sHnnoosZIQ4opImpLYvg+LIc2o+Ip6Xno7hkX/PGhMAcvzQOL
rU+Tu4/GRurVT/5Vdl5iyKsknNIDZCW4ebqaT/HPi8/GuRkgI+lKZODkzkZM
xRvwfLbsEFEZ1UCLfIhpEONvKzb8wdF0+e4aUhxNJE3A6LOb3Q7Uol1LJvdR
xWD+aRKaaP4O7TFPRX0wUXzayxGAWZhZ29GyPWACI5wb8bdKApkIPnxiHO2f
0i9k2vvDNGMJI7y8to77T2AoGy22fulQh2VrvSXJ7nyS7Q8WZM0NAyJa99yg
w8sYHe1Rq4P3dglKb+NoogJrzouDV3KrEDjNpqOcPky21jyNa7aRvB0wCPqR
UqKcCeL+LKVcv+SlYFbqsWTMc4oQJskXK5AUNX+j9Nm3DfTuO7F4/Cmu/e+e
XGhofzqFN5VbTGNfSW+c2lnv5bnfQZhmhgzIrQvlyllUMBUh+LX/ND7UncbA
qMDC2XMPjnIKvD8Rj+Pi3xKLSWOeJf7tlCyjMHOWFIfVMLXXgosandph5T8O
dvBM2zdhzwVG862H73MTPlxhJLICva6p3wj84yhATNY177vcIt7+KdqfmBrx
yJO9nvsHH7N97bjNZQXxCvQssVHPO8H1I2qzSr0HKNJSsGQo/xgnNKzfZEHA
NKkfLQMbu2n97TLd3Yx+mQO52OUGSGx1OeflDTCu81tnyDUJg4wYOvHVcZkR
zp3L8XFimDm8IlPWOcAfWx0jFBszNh/Es2vYyohnmXJgUC1fmd8WlD4E4OF5
OkaO0+Lvrsop3X4nFf+eBbYkYLZnmCE4W+pQpYw0dqa4MAkW0zshvm9N5zVc
ZqYSO4y6NlhqkxzVVVy2BE14+WE0eEDv3bxthaSVFcAByiZx/4iocAn3qVRY
aYf9oiapaYDSwtoKM8kKlsNzfViGiwCMeCV+C98lW7xqzRVg/Ajqt3iuva/f
qadgWkPMujcmf5B5OYHBbyZ/IeKDFr4ApftwJhjR26CxIlN+OTmFaXh0OHR4
8m1NXfKZ94BtLbk+zHKAWNOtP/bsABmRpREP+DVwmkD3V2PsF9PrmO7MRcUZ
Gz8mU3csoVGHA/oPL0eNpq9MmotylU00S0oHYdwPL1a81NRt/TOXrcCj98mI
uVa9+qda9nOL55QdHKfBa3m2rz5BStEDjlqPHjnjLrJbnk3Os63uLskjRpYk
xRRs8Kni0dg0N2r46xaB1XKy8+y+rwCf8oBkyCMIFnxtqSfo/Hbhjh8SNnk4
O7k+FXmNlMZYMNKPHeyFYVw35CVkFCrnS9i+pj6itMGUMfbmG8f1H1e425mJ
Txsi1vUORRNQ6zV5EQ5dJ3ORvR5d6uPTHVEAyTdmw/zgVDk83KebDjODhdqD
pePh/SNpSvtQWsi4RIPHwATSjMZUTFMys0uaryI5YmSWJb+SOw6U5S2xIbjT
j7Yc3oMEnzV0u4sIHGXsHKham8IE+laIRBqvLR+r9HuaN0SVFtiAfH6CI58Z
AGfJc3GkwcllRBqaOylVhxp9mIpe6Xz7py+udVx/6PI5wd9/rMET6jbIGFLc
MM2NFHn6J+T2z5qC8bydVFepsdvFyuKZpy5WHtLdf7GVvo44L5Hidhe8zSgZ
agUOt17Xdasls7zdR6OW1jq5cjQLWHdN5U2Syz0dKLKQNgie3933qhZTfxnp
tp7QDFJP+ZhwM7c+veT5y/+d2cFIvr/xBKXFHXCksSoZYg4LpO/FAiZ9u0nl
m16vb95iu/nh4uTv/en1ekbRz+IkQmlwTRpe8EWB/QJih7LaZmL3Wf/yXCr3
CG7mKiqihAR82taLz/ZDG9EBiD21M6G6W02TwoineOkmMtecYsRDYwilBMRL
53f0Gl309Uu3k/j6oZRoaeq7XYXyoTijaC6aWYaViw7PutCA2VHfiLgUM+kP
337AcN4JfFYUn/kh5x0SQOoKX+R4pxn5kI2oyy9aaoJdf32iLw2Z8L82umdW
/wXvVHZbp7w6/Ob3zcIxGGBlCAPmpMYWHeiWAI4Vs9E6o81w8/vtJUwBMqxO
+HZ+3ZNl3elnK2GVo9dsBLsX19EXlaT9GUo1N7uyBFjp1rUgWvKq60x113tv
5VikAmJPSikqfrBM1jwJ+nADUKxixUa5BqxzBje9R0CmRUxWi6QO7pFcPdvX
4BUl1iPV2Jfa/uGDejyA1iPcJEoYu9Dy4cLL+kUtEg9qxfD4kd1uyrYe5vzM
y6CU2Sbn77pGVfyVB+sAZGXuX0R2ltF3uufWOY5zdeOwU97H4U/JbYrWgw7y
i+8GkXf6UbpS9lZLzsIPmw4LC2scSQ6g2fbGk3vJ1uqondFmBQNT2M7TnPd2
ItaxulyO5Rn6d5JXzizQQLXOpxkgbcQRa59OrXzEvo4jj8gk/gEOyugkFgBy
5/nbejZA8Udx5L8RZMwJfuKSZ17zzruw6xieHI4YmyB436CRPg2fy7iOX34t
kffVZdM7aEthL1sDbYN2ALAG8j44Y8Qcpgi5GsP/n9R4pGC0Dasw/F7QNI14
8T45soR+trzVpXXY/jliZM3F6gd9nLozJx95TxhjuSKPV+bW9VIJCNas6Ri/
wP5EXBCuQTQ1RIyrD0/Sxk78htwjTFoVMN1PucaPpjfqD7TActANeTIiOylq
B4LW9lRvuCSjAHM5n2E/QeGdL7l5zvdf54kFsQaCNKHYLJWuidba9SDIl/F0
45A46CD+DI9USky7Pay0poafdB/qp6SnozF5xJE+9L7+TCYsQ4oO4vXP8AVW
TOaDdSOB4fTD22zEoawYa7qkHvsrvWdPPNS02NWbywZKw8odXvqaLy/RrCuV
LtnxkkbjEIUxOpQWWSFj972APjHZ7T7VZ4AjmNQ0rMJ3JeBh0ZAvLjarygS1
tqpWkOk9sdGCnHOkMo2A01s1++w13ZPWWWeIbxEgmRSJYLLQsO/sZquQbHVY
JDsaJC6UJtFNOvUwmIH4daSxuqRK0Xd1sw56Fcegc//+dJGyKaCkRhObj23h
75Vp8/NF+EH1GRIz01yL3BOVXysUGvSx/Q1YNeU05VE8kVTG5WNqBP/iXt7y
25NotP8f7F04TJeHUX4qNZWV9ZCPOhca6w4YlXBZ4ll/mW4RLvYrCgLq/qjs
+hkMB9kYDwO0xjEtoAdu5uBNOhsFsJoSNcgOFXVy4667HT8wznJR7cmOjSv4
AmGERrKsuNfmv6kIbuYGtUHqRfL3H0hu0xcL4b0+6x6phLN3WvsYPfKo5+q3
Jnj6d9gGyK0Xui+0myoKyvqF8Q733Cb0nrb48KXkehNl9xB3sPSnpDiNA5GN
dtMGDSxHLPAZGm3l8yGmlnT+f4XOOZ5RA9gy5ONStGXbYqlZpsjx3UQVTQaM
Hu4vRLjVGbh9yRCQjDVgBBmb1vQUbeMX16QRUZ5XbCfR5RNOL7KshxZofkbK
7udA66Xj/oRHAyJWSN/ycHfoIVTMzZ3oSSSLnUpdfHdut6UwX5KxDN+EIUin
BQbH5bvZwz94DWXqwVEvYWPYXq7YqS/cK1WXOQtCGQjAPO+V51FCAhTYt2aL
NnOVPDjXxIiC0sBuIFdNhnynvSQ8RnuiKyQSLWS74rznMZEtxlCcSiaOjLD2
ribdxlbhtrmG4zIC6GrdNb21LMNoSTGQ6Kxpp5kCvAYJvqchjQmKoKEzKHa0
/ro9wQHVl4zdTdIRA29N/1hlcdPlATvfsjS7vnIf42L1apu92Egl/M7R4+ss
pRtMLk+7q9HSeGb7OwtKihIZe7bGnKSOSgSf7sTezw/lcVJ/9BEZdSyvzLkQ
pxY6DIks4OGRwP2R5lnXxT9NRw1yK6gFks4/DANPpAdklPq6A3Ep6iUh6tYJ
PX5e4ZXlSkp4fv5YoN7DxuGwm79ovZI2hF2IB2njTItKMiWNHC8Znp52nPAI
A+38Pw9APswM7AcWO6k2Ld40tei2J+j1v6VotqRERpfaCMIpb2ESne9U/iWO
5f7eLsEjFUBcePkKyal2g7Qt+ZCIXxNbipri+hcVSPoxDAGEO7n3aU7ghhgJ
RMxh3xzyKdfR3lFboihr2623BKSDxh3MuoLenMAapnv8n7O7lQfBaZ6FB/bA
Trqf+eDlut+2AjrQokpIQr4OOyz5YzpBXrCyW8dbuN7TJ6tQnfu7/RSUS5ef
KTrwRl3OvGgAQ7229wgIVDvzElgv6o/wQhY/a0HzvRyyXXoh8nkhVWxQncZb
AF7oVyyvGDhcpx9vNsRf9ttx05546hhaZVlHcUjn8XLwN0jEWlc1k+MjSqNk
fdvb9JaQ8dMTWaw5fe7s5i4kWAeI8Tq5wlFfZCZi3aXrlwGu0sRzfGYurzXO
89EFIBWjzpP0oKVtRvt/tQyQNYGfTxehd5XWNdClb3gosUFjwISHFQEKAdEC
fj6K5cKjkSgJywJfu3c8b1JvVsoPvJOXbcrtLV3rnyu21bWyMTYZnvg4/xun
4cxUVg2GYtItuHDhNLik76lTRseURRhrLogMbovdTsowazM5hZxBatxd6239
s8jZZoeiPap8WMfUZuAgMKYVNoZdS4xd0UAg/U68hZY32QNRsClrj1YuHa/v
bXYiYvqybfsiH4xOtYRnjd2IdHXBGhsvSs6GlIVsIDNFkb+/UHV//VbZgmq+
RENjj3OJ3Cm2ajw9mNL+AOIiF9Qx8gfV0oo4OZgjTu7x7TO4Ivixz5OCLuDi
8RLEFVV5UnyT5f+IivsyYB1BdcepnCnBDpEPOWIO6C2RpkEsUVGdb9uwsNWn
tcGulezh3AK7IoFq+DhFYfD4d2VaI7eOWrByzmNAUbThkY3669gWDm3Hr/DL
eUtizvxjlmM70Vdax8kGeGTbiB7HorQ/T2BT8UJ4/85U83CxTFcz/05CoO9w
FALsH0sar5f+xgSsFy9vfo5XQzgsJ4asuCzOAr0pIvHFniSbcJMM/kQ5JtDg
ijnH+Lb8qp/jQbIUGuzVLOPQZWNpzUIuyLRhW/PNCW0eI3NaH+j3qSttj2Fb
ox0ershQ4cxhrOKlO4DHT7u7hhr2oOkIpuQbLb6CA5A+VsbR3G14TRPfH8mO
augYymvYMvOCGWibtZ45FTrs83aVWyomHtWyJYfZ42P5Uh/LMuzHwPZpao02
ZLxOtY+VxJ2r6/2/I++v4IjSSut6qrGaeKcivYEaw6vmgZo82edhJ6b4MYFX
AngH44b7BqkvlXxVVK6Lr4SplZOKcBjDMAfJOVMehi5hooDNAL1gq0PdFESy
a2fx39TOjmRq+wMtPs+yNYq9wwUaKZMHmFFcpyoJNecFbBCecCOw+mhxCCmr
qphQbUd1pn5wyO+1UGn7ILvXg4WuG0bk0hCCnY6Gxm3eaMVpDaG8xPe7YkC3
EuX/HuR0USW0Te1NcvByw2fiWthQhxpZaeVDBwSY1e4Idrjl6bfAihrxCZqM
XstPfhtRbIzdP8koVaDi3oKO2fxiKPp8NJpzL/E1GsgkQQ9nnrHRciQSu6Jf
XQ0iapQFMTBWk43fUu6k07nScXWxzOB9aQatpfLDKVIlgW8zLw/m1Bxyz4ie
vmhGYF/qq9mfvwEHUalnRrXpUDkGBEjTcuE7sZEzmlKlZ+6q8YvwiA8T/W7N
4yARAW+1mdCNiVX657WBvntom2FosmGwl2LN5xHCXskyXNoulTZ/I0SkCCsp
S4y6ce5ql7bPxFTTy2TsTux00065MmevUl/gkIZc9z3sccuKsHalHfeK2rjW
1PZXe3EF67IouqVcCmIgGB5BYYV38E/H0aEDQEsRkN4tcn6AVP5H/5LWUbKX
+OXnkf/WS5tVfRS2bR8x0r1tzGs1jAc7+lcwZFkNLSmx0i9fiaHu9zO5Abck
PlLHOeGj6ala7LS+3/yhLfvarse1Wy+E1quUnkRrEEDVAY42HmK58me/jjUv
CxgXHWVCTnp1g7T96Kv4vbAieUsuBUjob3yoTHUSYg27sBr1ANtdKROzOWb0
Ycu+fXARJdjPzkwZammn2Fo0/rMrRSAnIds9gl4KQzMEZw+52Fk3W9uQhHPo
vwFLk04t2KqRDjeH+UNr20UfBByK5AyK9o2gnqtQMfKJneQwYLRGeUWCr/Vp
hz+KUGX21rR5UDl7VegvAszOEfYr27YFcvsBDYjEGTSRkNw/M5sk9QGg4DSb
B6wJEpbbRpTss6ZjBzvdaxJyVBYaF9ghB6NtGhAMvhCapy/pOnjvzLdRlYqA
pxgQq/IdB4ENtEhpAHE3p0TOvo8MGluCfU75iHNfct9MSumIe+sV7ay1CicL
TYazjT68whOVnLh+pB5gTfeAk9QKifYzD8Ip/7n9wnCJwiiase/r9W8bsjr9
WBUnltXz4jdvh7Z2vb+O/MsaNnPQ+LHSJ+ndEM4ORLcT1U1nioGn0X+Q36HH
tCMDF/qIU62Gd0AZFbQ/AXLQ5CrSj5voIJuDPflqwRSYnOEd60EmHIoWTBfW
Aj41XwKPycxIXCdb/oxzUPtq147d2mYr29KMBiSaF/pNEiNt9Bbwu+4ef+Ek
NuaLEfH5Aq0n01eXB6cJ8uMSraQdvRut6ANVH4L7cEvq0r0NauE3Mi3XtsRg
hp5wMh7FD+ELmqbYBhIHranQ/gpNxIVCfcwhpX6Q8NEk/twrWkWSototDyBq
ixnfgDxO+079wYD5m2b5j+74PZHjX6puLezruQ5RKsSeMAzhFnITKGcQvEw4
aPm1PCOVNvGHBaD5KYhW7RlaOKfFbEXDCDu6UjPSxAC/AD0LLzu31GhFrFOL
or/nAw7UX0b+58tPSEsxTNlBUxsRIwY8ZYBUk9NWQc3JIf9QDOhkWxwGQGet
XrcROxlqEXnvE28TgCMVNg6kPhp4pzEiMChgde18jEV6cjbmel3/tMKCP68g
/jg3yC5dJrqACrXuts+TE448peuaO8Pa693+8CctgnPNrk4A48MzF44OP3+V
X0KD+u7+LoTmvsDanfxaLxcAbI4/wcu3elQkQwcdYepDRSvX/XX4LuHmalPa
Rx/CA+Kp/VvYRCmoSv+Qa8i8cRNaFiNNb5u9iAuJoFMF/gN4CCrGjKXJerAt
2eE2F5dWoaa1xFb5NrcXbfA4Kqzyut0eTnWrlicYu6QIVmwUrmhuLF21I7B9
IN/T3TG3fB7AE8/CMm90W5yt3UzScBglj6ngpmxhQKvmwleV4deP43dAVxAL
45vJ3u0CuqQKWxpM4tgcujbrLuhiCW2wt/ysua4wJGHaS8zddqmn7U6yOfbB
IuNF9EDQnYal3CBqg8mbbKqdPNNJsqpCA3XtnATGkEo9lTTn5Lyhk8pKQrxI
u6Vz6zLS+orPZHw7u0IBdLEpoRP6zy3ZzUvR+W5I4o8/94LM+ecbGyWFVx1+
nEAoxz+Hg9x6KA3k3DhONUGp5uYF2KqfipYkxMoKAJks3oWj+c4OkKESvh6Q
gYgpAoSwcqK0iQtFivp6Fp/8/B5AYymxNbF1PNMbZlBNYf3SFMu2E4INUNkK
FB59vBlYQbUTYF7uyLqcjbu09vSed8s4uAEdaadI11agegjUg/nvhmcGjCIr
oUdb7G54U3rKRJ6437FoEtlisM5CKQMb/spWpv1Wm9KotgSD26+6MBxFnrMV
BNd31P13XqvqCmzeDUqToW1Trpr+8ND+DPqT1L91lCP3/taO3GGXPbZYarXP
Z5YpVUeZyHYa5vP/sjOBIPslbCW4qdSrrsHqKv609ssCTLPmtQzIjdun62P/
wtmhP1rbqGHWaCVzLwwby/yzrIVNMbO4+7X6cl274cM9tA67shODVyJLU7Jo
n0XJCkUzq0XZVQG+tsih2jxHB3BQxOuR0i9FgJZhXr35JIr5uz8s0cOUBC1J
3JHe3ooQtILjczy9i7QUgmIIdewhX8TnCJx8iDdVfNNBcMpTCyLlxRCjmJ+y
tHdy543rSteR8rM337boSXsRG4M5JYjtXXN9C99I/vlL48+1NBBvw1ZZtx5f
mjshmnBqu4qY9U0Icn3J/ihAyP4FydP7uSsVc73JE3ljuqsckPdw8X2A7QQ5
biMJ/NjuyjJh0j3yhORgPLMUmnamn8+cOEAJpJeXbVTRe0LrSjwFJ6jkCkKH
hoFs09l5wsVAe84PISWOzwHcxEuMmLTJ0vzKAzeXNMBWbBqh43rS6+e6tXVQ
oI0seikYHTdYM/7N0F5oTdfrJ5mBXyCmHGHVUcx3gGWzX7mh3gtPzK/uPU77
1QwwDa6KNWqoF9umegAsyu7HsjPndXq9rm3GXnPdvlM/XHiNIl8WufpbS90c
u3Ac6mu99io2moE+xIJC0IIMaKgh9ZaEJ849toySVPvbTQp+qWbDNZLeMypO
D3E9doPLv/jdmHtayS3emgURkBl3iixWAyPnw7+c0qRL9lD8myxmNXOpV7Nr
nUfsODqswi8P3L/56i1Hl2L49RV3VU8BQ0F9BQWaQrBjoTVU+IoQvXTe/Vqg
Ix8MoBPfygS4NdVIGDV+VxzMOBxGsmwtV33pMa41BkkL+gakJNF4sIwlXij/
LrzY6udlIG6FevFqcPJ1X7jBgVFmRdlGXizPfAltyLysHRlVzyzdBY/hrwHE
o/wnJwW+fPVejmT0gCJxFIUZ85nNjRJlh4M2m9DrPmU8rXm6ICy58+mqA2rN
1MNud9l8dm6/8lzYCkCr2ODeVlIjNjL8nC1JKdlOdaJnr6ndPEIwVn7ezDb5
q51fw//4ZMKCYZOpK/uE3kCTnjnxWI2uzgh3UUzqkJ/tpAurk8CutAvlh8yE
7npX4YoUxfyi8dHqXuEj4+GY1ZSSdO40DGWdGzb+rOhHls1eWtWUQldfS+ye
x6eTr2NmPaaA2CWj0JCKZr2fLZQKX89+FoJgKyzBdP9fNi1ZDb3c/73XyaI7
KJd4EgI1EYCnXK+aCza7Heh6eTFeq5fblaz8a4UV7++dA2q2d6fNPprfZ1gY
Jhm/bgcaDjYFTq9Dmc6G4oAXbnqJGxsfk9ZO/m5PQxTwPMTCZInKA7aeMbKj
4UPRdQggvISMlFdBKnhM32yT3BTeMh1k1LQ9Wd6d7Djcvp/7EvokGHZtYMjZ
toZ9fHnFdx/1GBTHyJL53Jn5s+bNEy/bRzbYO7oGRu3auDbeRm+r1i7yhNTv
1LKVHxktdPN34py/+HuRqNqEfKyC981GyPQkqk1aPEfDj/jBe8JETR0ldpKd
Uq6vkOQXQKXViIV6ePbqiCw822I2AFuIcanfvmUGdttceGek0BDdopJIR6aH
bRS6Px2we0ttz/AiFXjhgq3h4xCW2HuxFRYC723cyz4xFZA2G+0NTCMLDt2S
FTEfLdAVwl+Y3kvEUrgf5SBYIOZEC0OKl056clL+/KbZJs2mfRqGJFXQeQo9
KVBWFPD01d7sw20WqWdskC9ZjlwubuKP+IX4ViseGDGh6usMxolgxhpF1lY7
0oXZkLI/BXE9R6Eq9WY8PDO+uEVTDDKL3kfPDUHgCxw0S1YyB0eVAg4ruBTp
DkWFefr8ReRMn2jIf2nFpYknLF+9ivsXWEgPxAQrmtOdLAh2qJPmZ9FlnrkV
BbXjx//QgRzUuIgea3vX808AUtxc3nYi1Xl8YnEsZg8fkEFkHjW46C1U92xX
c/1o0mrEEgIu+ca3L3GBoWsVGrk3jzLRLvGgoSGsUlFH+8PYU3l0AeCChp6A
iIZCNH0kX1COkoXa1kwoPxxYxAXXiX+yWhTu/PDx7AJ5Ru+yODnAmKoQh10c
xLMmwH/5N6wqWblxFnub3fGtMFWrobJ6llc1u8vN8G0sAUTSKf1hqljA2lQu
srPxIwoscVCiFM50ha2aBa2zAgPSx+e/ZSd6AhFlmwG/nAQ/9YfvYMc8R4a2
8Jo899bleFoqpT50PDMkVTkoEwHpD1eLBEX4hCmNNcPp2DKfcvvyaXIhPUIi
IFDNHxfe501ocmhmqKzWI14pnMn9iPlGNq9J5IhKFurCIrN/72P7XbmMi4DE
JQXsw8IpxiywRqKV0+ktuwS17Bg1LbfkylP1cEkq2JfxCM4zkV2YSAIbM6Ol
a1i9IKeBxp85Q5kgoVLZsdNnOpC7MmXaMCs5G/ZGroKhhbim+Vv1+usGggna
r8lE0XGkpl3Qx2240lbBbJBgMwvnK24BCxpQ0X8567gbVEHHk4HIrb+D8Ar/
xrj9NpA4TGe3RGN0ch4XtTWxuSBOm8J2Bv/yP827vkT8jSJLqJuEMRLui6bf
o/UjFQ+ymJDGLNm/7afJU1Oj0T7xNSsYT/EI7W7Dth0abQUX0XPPYWYHMevW
Kvjk/n9NIeF4aSEgTg5/TeQIS3HEKNKeWY+K9pNsb2keOTMm4/9mrIwolbR5
ucS3uX9sSTt4Oc8Ioiw/dkSp0gWjINLOkNXp5Odg8daQRVGSpA4ZUaJGV346
PCF5n2zgZD1nLSzmiBCHADJHjaT8vuQo74JU6HanzASPc9eXeBhSjsuOueaO
qPFTJhVQ/o11JnDpNWdyqs8yL8h242IP5y/HBupPDc8BKG7GGyJZMindNUYQ
9f2OF9Q0xwuDZsYSyf3x/bNhbrxijkEQ+hbzljTlR+6yXbs9ob5QHCjCJjRF
mg+iZYkjhsjlkP0YooiQdwRetihGwHVb4AHw7xx9eDWm6iRa80oWs+tJxjAt
HMSByELawPFvDoyh68d0orbAMBiZCBKT3nV9McGfeDnbNNdgxp/IilvOleZG
JlO4+E7DDUgmgrI10kslCuFEkwF/RgtampdSkskFPuuHsoguGcUkr8FBwAWV
g1WnphY7E8guzk0M1Pp7YOGBEc1cBPxXWncsg09pybpbYfIHV6yowctWYBdy
b7lWGrMFXBOp4AGGMrkTDstdpzaO2IEqHzkI0J1YKhW0sghSKj8ytJizYmRf
N1qkOzyRHfcAzTUE3BxRamknf+ZrUPKbaEAyFFobThoxD3+gPtj/ePm2YyBK
LPZOz9HJFNmW12/AYGk5ZXbbAlD9hFARs2GTcDEOdr6zO1X9q96IxgY8lu0h
3wrxAsoua5AmwiUl+0l3Qo5upLhCJkDbmcfo/iumT5Mrq82yhD2oPWgcXM4S
DloSXDPEGqfm4HD3Wxls+r+z3iEYljgo9CGJvdalmcIvxEj6rhXl3xNlbTs2
Idscqd6z08fRTmV0++BX4sam6Oo/B2CpZhsv5To83YJ2ZPk6sOfDdLeovyhj
UW0Boe/a20vbpQCFptpsx7fngGlp46R1ni9vv7hrHY1/AWaeYIhTm3u8KDnj
plZegf4kwoV9mbbho08pbzlM3peHUrb9cJV5uDSzwjjwkzqjDAYb6wyGY3vd
myT8ljyWvMLV9UnJNOwMm4hdiKFiBObnZjFpAOqTAFD55dpysO1lE7u/k4nh
hHviiHNcRq8L0bBSGRsEj0u5ixj51sbFYW8aJEiDyB4uCHCkSGSQfVp72cks
4/oYhGTetCbPYJyeKt2eplLqZwT10ZKNBTLyeGciXV+Y7JOrYa+9PIeo/HOh
P8qdiyLfJ8RK9rZUnHWQFzbU5Zk3X681n1GKKr0NuLHp00vJj+QJdfdkeGO4
T17J4frayFdpbEtD0BZk0IHWl+eIu/gWt3zFyxpcCckU5h8oYW309rJxVsi9
2+CXLZujvsHFZy0eYsQEnU7qJ7frZIg+m7mBb9R0HkUZxgTscsRDbgjXrUVB
GCZCT/8cUoY78PEMZ6FTS8/2ixeu0WxXd57TT5KjPgG8jrGMBUHiYF2yc7VN
302tTOPIryDYdS4dcZWwXD/Y5Pn6gjicLjSk+83micnyVvTZEKup+T+g0ZQd
Wxafm+Z87582w6NPCBkwepiUiOk7lr6skuYyt39Q/2McFrJ1z3As8jLD7HJs
xLHkg64EXTmZaxltMhjxYuZ8TQVSltC6uB7NorhWVy+EawPvteiqF/lS+fes
cPe/DZAl+wW+GlHxSzCaQShuVqASnLwk4ZIHlI9LQ2dbjeHW6hdFgYClzGSn
AqVCNU909rjWzAq6/obq9twjRKNX257RXKQhq5BCD4CxnDG5tp4Lzo7K5ovY
kD5DJhzQ1b+dqoOg+qpl01xzTUNWfNjtHbmhJ0ZGUcawYo6Vqp2cLFdLYJ5V
BDpwLYs7JtjoIOBnpxm+FsANYlx5Iih2toLzYEN1S/ZVRiXlColVuiMYv8XA
8cfontH1U/sKyUMrbYyRpIL0NdcLIFx24mZpBZ2F8WjRdqP8fYZ1bpDVw4UY
V/xp8hlmGTJQfHFhJ8gmpTEy0lAzYisVOMXDOciPMzC7lqPxSIcS20Ea4qzl
H2U3iSKDDb2JM+0gpM6uF1E3JaAx8tfyR9gLFffsAq4801eqg+lVV/kUCF3n
frO08yC6qechAYie0WJ8EjBEyh+pLrJOA3LY2t1nQsYvqoPqhv/z26j+9yem
mc7u8uZLuJjrWPlRGggvKZfF/zGFzlcgb+gH+bQoiOg+nf8rMCMTIr7/RBYA
WB0dO8HV3c5UE3rxnAwPd+Mk7aJJaU3hCHVbV/4ctE9lSRRk9kEA5DbeHwRV
sJGbov6Gx+1D5U+cm6nPd4cRnAdHiWIoyC8emHpHfmm/Cby+LG2vJOPFbD/s
sagZFe4tQ5XxedhpALEqGjIA215SRoYfDLFeSt97O39w4CMVvp2DWOuE252G
zYyiah5LPN0tD+tsYEIAUuKAvB04v4y/dyAQ1mjaXNnDk9UsATaD7UWbA0rL
GCGQpe98+rRISf1vNwOOf1YlSE/Ws9WnaR0NnZAAIGW8kWDMz57rKH0pqZS9
lwEqZDFKXkQ88FG2Dmdl9S0/jGT6D1UH/UyyItYarX+7ZklwUhGllnENFlTg
SPRz97XnM4dNwRVgHmXiBM3cwcO5L1svdB7aUanPdG4uXehxpnxD5SFSZ76N
yeX9nIRJ4y1nSov57VCSvMLJE2LmroJdC1TmPbrLV8QXS5Db2qRB/Q1+EonA
eZJZSc7AL/yHJCctg3ZuI66fv93CexeTDoHDfCZ2zgL9fpdGO3pM4+0xWtQI
7Htosju6Pn4x65abIfLCJOTAZ6RNvHFnv+MWnTfMzY85ejxLZtRYT72Zsd4D
69k9KLEi3y20SoBWeYL9l+a7eYSRN+OS1PnrFSEhxWsWfErYywiIYbhJeTU6
OSZsBwOpD76XqTV94XxZWPZst2G7EQuMkqnLbnEObhDcpFI+QfQHkdLWs5xw
a0ikEVYsMKmvu7A1/KuosNk6PivbTyIUqPePVa3UlqTdea/kODImWTfLYfLp
i42oyXypCOj/dXs67Ch7cqssRwWQkjYLdZhm2+Bihen2DuI1//mzgJkrCJZp
OTKW4qLIZCelCkffJCtDbxbzRMaTp9ovYw7p8ScacriqRTjHTweHjr8RMg7r
+zcbh8EJsyjlzX77xEfMO4xaF1+5ufMS5nOOkQ1tPoWp7P1kokXYCFbSmHz2
+lSJeuIvqcmnzwiQZr7teKWVOhbfTi+pcxn9U2nIVNERwMV6VH+or7W5RGHs
pwA2BKB+JZ2i1+DyL3lXZH5vyFNKzMMNkgymQN/1pxRHi1j+ejS4bVdxyg0A
ucIFhBWFugi8StNfopkEHX+1JltOzL1fIimMj+SDy410lLnEAuIgSI1fhqo7
LIFI50lzehjTcIDjMSQar+drS4qEWYyvD84001PVimuLIDx3xM2GxORfmBbR
IDpD5kfGARlJH5UxKWwXtDEyceoGAPdGG5pcLgpzQls0GLpFMpQ0w4Z9GTzA
T365IvJAhR6o+QgQZuwmAHE7cxm7NilNZ0cMeWwz3yJsVGRdfTOhNbV/n+0r
iovckeflFc8pk3+oMuWC9BhlJDJfklqt117i9MRqgAFjnaxqJyMuHyb+LWK2
YDakHp9zw2654LSINFOyQwLKDyJczqhPGzDD/c5CYQcBRUxaPipLtmeYcY3G
JY6J6PMtEysq6EYiarIeb3yVV4BUObOWeEj2CZ0Dm4wwuPnGkv8+G+KIzopi
TSKF206oPyzHq8vDntOwncu7RESYEonakxRHeW5qm2M67Rilm8cIETmKMbDC
ot+Hzs56MxikCrP44Fiqsvt6ZgWtSbnUnXdq29KQzDc1vkmZf9GSunmTuJmd
gQyvnjE0ZtuG7D4UagMXtM4jex5bHRXocHymXtAjQFyfmDwkpKW3OMGpukZQ
49muSQw5LIWu+JZZI3kv9F0b2cacBouwS45nmYwDdhE/XYAU0QRzcdegKPfX
XlNmnX7eNSLYb2NA+TPXxjTlvygoHIkjZYDq+UpC5gYKunIE5C5ulYNegfxa
K2KH7Kj3VCiXKUDO0zHVGaF6QGJhGXjTGgrOEesdv7VWn9cde6xDoyrDPf+E
tiG8fTOeQk/34sDENH6riVqVBl7+mhNjWrzS9LwDvj9PNq3gavuSRnHGaoRS
4KX4+SfmkA6NtcH2cqORL9DgV11/RxmqNjPqRhX7tyAo1NVAYeyIfzwZIS1x
L1Nxuu+l+xYkXUQQ6jPR11TR5Qbthr0z1Aflil2FN5OLDx+o6uNguRFLWcZW
GgrIsQ65O+gqN7RecXK69IQvTKtdDfXszzq7vWBxj/FemQKcN1nKCo11/8/f
pKMdsshRmWF04p6/NtQ51uXNd3KGqy00kT91PB2JXAO9mcmpUiUnOPSpKC0S
AYctdbDp9yOIUpCpmot3U5p4QcLLWOM60aPF+ytHN2/3EXkmUyd0OWZj58SR
m3+5s/6dpNBmmHEUalk3laldy+MMXzPuzifzeyidl6NEB+PUpPARElJh6lIN
EEHAEoxeox/nMLxezwEwsEUyYJrxRQ+oCBTJn6X5Yt0tF6MtwSpJ1jF2Ts3u
FsnPp0ucTG2w5ubMUND5au1aYQU/qGvgBp0RI79qcce3nNpHGrDR8FqZTitl
90WgNtT7FIkpyQxeUzuJTIHWuEz44Ji5xCjdqlnmcv6Rnx+E7+bKTuYI4IP6
ZDZqQQ05xizTWzFxGQsrLxFkks5RYQPc9YIf0MHPZK6rJP8GB7TqKAzI3gxp
DTuvpKNfxUahh4Uf6845fdkugoDbqF9oNk9AZGnReqxAU6X9T01TVyDipZBS
W/vsMaGD9URGSpVLF5BV7KDj7CMtKimNwfJoAAhYOxfuANbA+uveHdq+qUKZ
GmgbDqw5TFqsTlRAaSIfVQD4EwiLh0YBVVzxskfiqAunKnImp7ceNorF/P6m
aime3jqr+pDDLyY68RYCDowUkueXVOnlEHUwEGb72b58223+QaQQQRI56zY9
dRvib1KWUxxtRWT2wpr9eqRUAWW78dt3iL3u0tS4VE22aT7fhlF2pJbIrlOt
gbrTeXnsrwWIBgZl5zCSPF2vR8VuPPFKHuc78RikEH74gk/dt8dFuf2z+6Hn
fny2U2PGY8Cn/zhXX5DZnZBD5zEuJZlgjwDzlqGu9f8vMExhyiDLM7hRyO4f
Jg9ubaWsB/rwrWhMZnZnOhkpMORsKevaOQsOT0YOsFK49k9ap2O3JRkIGPaH
m1Fky2VFAhoRRVv5mW7WE0QQFtSudtxq5aH6eZOl3tVbCA8pI2nI+JdjqDqX
j12IXXCQYpL9OVmMQaruLHTJpIaGoOaXh8RTF5LbdJ6tvDYmGj1p9igVYdyx
hwISdXFM4HybT7pIoAaqWhyJS8iR6pZltH1xvWvsUfDzEhwnFcj9ZIdadHee
z4eNSRFmIfU+mGbIVBo7cqyTkQlMY6P6AmqEasRI/Kt5s7Y5hpx8tHJ9ZqzP
Ei5V7hy5tpQa0ANcCBB9yfFKN+zo7HUhQkUXMNGvmCox7XiFrWGUBeusV4NH
k/cm5qPiAacXsp/8LVWjtNLfPI/m7BKEhgmqF/4EES7lyOyk3QKu0+O1T1+Y
m2y7EdTqZ5JUie5c4nMPIBZttf1fF1afgEcB9BGQdwn6vQwrJ/F3OpQnCXtk
FbmjAuVrtSgFsyDEQ3rH2iaTFPNEGn4NF2Cv2NtIftkLuKQlAdTaF+QCYPPl
6Nb8Jld5VTPkw/yys4S3BA2eJ/GNdb921emN2188entU2rRCNqLX9xMeFKzj
XA0qoiUvAScprv2KG2fGxBIAXE2Xm32LfXdiWpBAyugIIeLMshelJlId0hC4
yvYPVWkq9FSBftvlNkJ48UiEKug5iqKx/GaQSs/lNy8saBPyXFR4jOZrtFnS
p7mvKglUQwzrw19oEp+iWHMAhPqlRdxV0x0Z2nS1f/obYHVXF999ab6Oiye2
DLUrDzho4IuAwqdp0LifypSQBeMazVx4Tij/fONtoqTYy8m3uCwHUwFGpxzF
KVQXxpM1aS06iwy01qhXy0V/2jz3sFi3+jwlzviGL2BHaPrgngBJ9AbDs/CJ
feEYTmaofd3V2g2TfRd2G7aiaF3mtSYt9pSbOX+ROkkj+LP2m2l8djKyg77B
+QfqnCZ46ZnaXPaUyeR5B3j9BnkXLMMGsXDUNzRmbVSWH2UBuKB2MgqwPIYU
gOjkcP1/49vZ3rMPRsFK1iAgP8G2353jDBnMFNQ+biEk95luCRzMKhwEDc7y
EjUCjkM5L3O0EPGevskRnjheRSzIv7GAQeJvBdPa86CN8J3hvba0LTeuysuE
1vFuSUR5VJXWWGe11LfiNmtM1PaNrk8EY4g88i5/H8z224c8UR+UO2GSRKat
z7z55tsZGMaqKIOVD5mD3zYmPime4HTicWW3WGjKvu77/7LFU1C3Jsud2DP2
w41hjzb/d918+eEHZdBdFEaWbQIxZsxfdgDM8tFcqO2j+6NkAQkABmm0QzUX
578uTVb00lDJ8F4VWSdT2C5cWNLP+F3D9JsOJKWL9C9HB3cqnCN5gL0IiJiz
ZAhgCChrLYm1AdnrThmuHUwAEq+knkpz+pNW4+n7/oI1GjO0Zcfjx7QGEfUx
AsX24G6/FZhfT8mdPScO1DUAg4weMPr4qMcgBf6Rjy99K1osVt/F8ErX2pHI
gaqzyz1vlV9Z7SlNggoIzvlVXggI5vCPViwTFpBJ0uBwXIs781CqcKN6XHk9
6xCOKvKHx4O7T2KvAk16S3Bh22xXyzAWh7r+Bv1oVQ4aTuyNunmQ5JkCNWyY
5/rf5/nU4cFzumGYdBA1gRr67O3xm7jvNkRg3zhAUoTsIvqDy/N6zClXb+Op
t+JP6nqgJQ8gBcpjqbRF+XEUgf5KlFc5eilGKAx8B3yShC52uQlFk0DoPkn2
bH0U6a3F8Lf7jfxfJ707K8LGkH75k+eZrQqMUmXWSLTU9/fPnankZ8IZ0ynd
stTO/2+Jnxnx/ZWhGcUlcFuLyJqeJ2jtjOyQHJDsicdbXwbfoRdkPzVFrLet
4UJmEp4y9BawWCN+tTRyAQFuaaE5Jk4nUDPvDRYuK4prAjy2uGh5luS9DV/i
wdAmVXPibHqPj0+Zu+wgkFtkXwmcDkjGVNcJRsYI9tHNrjsT+XXCWxVuf7kw
r9EUkoNfSQSNipJpqP/xnLhclcyVNCQPNZBQtD2rol43n5wGUtOwvTZ+tfSR
V1yX6pjXlHph46x0cSVyKSYd81ONbnPCy5W2XL6ZaepFWlEuiGu8xMzu8ExG
Ar+j8CwJRMjRzJ1GWXH4gJgg1dE1uJPGIRFS24ySLjdPQOegyAxbZ0fbdMmh
P+TeLwpDZ+Em8b2nlmhs349Wied/MWLpRqQfOAXBfpyGGBnP7zLeM/EnthgI
Sb5QK9/eNv8LUBQ6bezm0Qdc47l9zkSA4LegFTLUE6tqUtXjwfkXBWX4uS4e
Jh+OXSGCNdK9oP7GE2V2Sm8D0RtupR/vYCDVkqRJXVZ058uvlTVBUaggx2+J
h2KLgMfNkcOgRjORQgysclm19PqT/W/IgvByLbXwBo0VXJkK821rX8RpWwUg
jSVKK6FpBQO+ravnfdtxhnToVdpW/rhf5rNN2kqvaJ73LphPHcVLKQHWs2F4
2gD2yVbfCPwo/8bgdCseQkU3nJP3vlZ48Wa7Jz3SaTnhMTOGiATWEmpQOzHz
8lOlHhxQC4n9aXs9NpsgeQAUABxpqBFOIOpZmSRQf+QSg3/0zATl/iWA/JVZ
OUKvn11FN+0JzDh1JIDTafMUJudPto63RaapqWoyda/ToRR3S0A8/KNtcjLQ
5ur3L9yiujcN8izCpqSE1/wm9QHnoHabhxDtGd0IGAM1F5QQZSokjuN/c3Hv
CCeEbZ1CGTOh1OFC7IAvi95fIZGpAjslRqHMc/ySsH4kSiXfub/ovugNUEc2
5/iVJHeHTQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "OJXsOzX3SCOyhcBXS9yryN9cWQxQkhDHUr4mzQikLKNKnB6JkSYY9xNnmYkvVOJ5f3SnsxLM71tWjwpqmyTCVkTt4jikDmXDCnl6lQn2TVy78ivgbebFE/F7GUr3Z8AASPmtz4v12cD/Cz7nTJMTG81IGzEoV1S4KsV3MBcbB+1TqTshtjzQ4oMMPpNw9ltjOjjqx8CktvtqLiQWjnKfQh8i3R/5yQlzObBDq+VCqANNLj0J6Lcvo9p+Pxo6YhOVAcwJNDfg/Kat+Lvcwm9yQ+9Qr2+pctX+eaK7fYDGfFGsXtG0d6mfND539NMfkfh9LizKuZbqoKmR7y8Itf283GKkDG9xA+NP7BPAz2CPGwiE+KVQfpiNNRhP8NrYU7hU4D3CHfysJKPw11C2qryYTRu0HycCe9S5J+qgZ+SJWeYAhj+LZOSu4JANKPnXlvwgmLU3SwzLD5j3l1ppzUHuRNN1m/n9EFniF4iIOWwvldI9x2sIX4yK1o59yORigb6d44p/li9Ll5JTqOxyEKg6gbRjbccH9KkbsFeFjY+YOYJth9WmHQoq4TZ0kIP6N/4+NyED/sSzO4ZY3X+RUELG32zdsIpEyE2fA1hh33nEHlUA0eaO8lKC2feqZDffiyo72g2lEzLTw8Bc+R+l6lRndbfDzUl+uJjigBA0ZkfE45gd9ju+WrBv9TtmxArvwMEP1J8fTu7Cc1x9xpzOtoC7kVFgy7YSU4Midx8nbrUqy5dbh68XSDlKkBlWiB1Hx40Wea3/NUEKdR77eC1Lh8R8H6CbWkp/SCckG7/uoYfPhpMMb9UGBPtMslMsJ/JlMYkLhZQd12WxNQtZm8sAKPwELul3xkHmYWjVPsYPEcLejb4dArZjgODpGiWL5MCBbql/kU+/OdXKH0Cgot5mSf5EsPhcDsVuu1mZBrgiFQLeP1yCIfdEZEWN0dGQeGJKfxzRgFBsgrm28YiK25LIZl/tuwv4pIuj/beQsHtpIY8vF0pY+eZNKRx/huLf4vP58jVV"
`endif