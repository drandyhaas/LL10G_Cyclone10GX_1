// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p6+BArD/Eyzh8EfO5Ue3yh4Zpcr9w+29Om+njD3YDWmOm9ZOi6v6vvALt0Bg
MLsugqUSI1DumNwB8Mxqc+vyiP6Gfa6LzEWxjyKwjlYKAzwC+WoZdgpn+Cyz
tx/3MYspM/8syZ3fOb3hvAz+0VO4DVtfijwnp2tnl3zk6cwQadwRrbO3DcNJ
7crq8zKT9dGE0Wp0ESETVTT5ENeu2/MnJNKDiUCUZL6RaL/0RxerSi4Y5ll5
Kj70aV/R0AoSt2M+b+TQ8mxUqBpjbx7KkzWtCKUoCU5bhweYIDGaK/GWMg0x
0GIdstJZkmy+RKnhUydH/ygv/YDheyYbc9Vjj9et+w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hGJ3e60m4r5xH/hueg4399sZ4drK4QRqBEKlKM45J9AEeeIoTOgIcGWchxB1
U6r8Vm0Q5tcgGkGrghevqGC2Lxh021Phqtzl2VGT9CZm1gJOcf+d4hQ2RGgN
rTabowC0x0DPrWFQCTgz+HZkxFOSO5DuXbT+VMerARu68kCgv3dGkUWnEQnw
fghnOGCmuljpXG7RfWxH/pqz3vV7ip3QJ0APBgsttzNqmcU+4aMKnRx0SUQ1
CZiy56g35u/MrfixtNnTzsGKb/FC0FDCpAd0N8I7IweXGox7tq5QCWWLIHit
bSFpxpv8/YQdWCoOrytHj4WtO2eiC8BINDw1Zu/Hog==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R8e2HYZJtk/bYPZZCfAQoF7s70XVeevOLtjpproRtC8VL9XqTPsPCCTSDev5
Gfi80Oc5ME5dXLod+hvCxhJZgzdgbWUTvmo5aLSsH/6apuVPMbo3YCecQQxu
rWxGK4JvUjfPCR71NxxSlaJ7yumFtKqXMyL2zNDcCU00yOSqOiLwoP7LqNs1
zPp/1Iztqy0hnfSucRBw4IqYBVUudUDaYeLqq6zSTZOtTIAANgQcS/n/DLsX
BMfOSY1BGSYlrZuLwppWvgXqAj0rkjCPrpeYU8hWI6gGzyxVBJjc323JEQDa
IIWGByVzkUfIjz2B/vjBUf2v7UXPvUgwM8Q810e9IQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IXmlbfs1E0mJB483lMgRyMGZzubhlhRUjB2/hTdWnCOe3dwvcp8vC1v6ZR1V
2HAKPQDEkSRdWZG7N6VWnBc2JM+ocnGTh113lWDYeh7ARsikLelAJ3PkaxiO
qKZMBB8cwi47LlekKcWpzCU3QK26P66r4x65QUHtjZtohF0/jcg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
OCSmPzFPZyU0ni4vlLPL3FnYAkSqd5RWZBcBtcdmIrDCBYMiNihQdf1Xd1PQ
HpQxSSl6prP7MfG0Z04wnBhlxLxNCYYGWe7XzOW5CV1EkJBMYpBMTO0PiHwv
TYt6ZFRNTJNAku2DYOjuFGNO8HOgembj9XfZ/99y/utMCVTMBpZtiMm9UKSs
DxbzFLyXjky1ialkzHM4YK+l7RSVlLrtHPjzgflopMYpcQuiC1P+gBC/hoxu
DDmMuE30wxN0GrK7XhvYC02kHq+39pABbQhzVN5q/jMB/5IcrkzK4AB/dmKT
a+0j1MowKQ03UJA9i7uqv0ovLmZI/1AfDi5yLurDGGj4phErCQg1PGVAOwy8
g9nRHYj5u6MGR8QAa2V/LY+X3CEldYidjOfPcXsnwg/+Z0+eq7ySnZy0uSIB
bVS5Q1b/ZyaAKMGUPoC1OTlJ4eq/aEJtNmJqTaaA7atXB8u/XdGKBGhnjiT+
rjfVz2yKKRW4NrvZ0x1fOKvGaJN4a+5B


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PR7HzHKV0S7QTjtf0Rz5ofJ/lxTIGq4hK6tBTaZ/UjDEcGj6x10jsClRlEgB
NN3mnjtD7wt8VHjtGLcD5OWtnyYlOTawB8qGEU9ULRDRxhTlCLm+wGcoTQug
J1+fJ61W8YK32CN/H8LVj1KYbYhj2hkBBbEUXSIlHHHRqB4l/Vc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ewc0zLo5j4gY5UOOWP+HGMg5qbGffaEvUIqnfZKMBwzRxEQDkHXwDhS657Z0
JG8IyvLbcvDKKfCQeA3PwaVEWbnPF1Lh0PqjKi1cR5Df7Dpdc5iOjXFv65fC
itX9QrJ5dLOP08DwPJGxuf+qJR60YacU+waz47dVQdWMGwIv/60=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 17168)
`pragma protect data_block
hFcqueXpcH1NEXxcAUG1W5d0O2Fxplvi2amWK1vNYAyBlgnOnbm+awPQx7N3
kZEjXUjJ8TtdIXw6ItVMpxd5g5Zy9xEjVD4A3Q9CEG1ecA4IxGlbrK6nH7Dc
PeZopIzjBrJRsvyQTMA6pjVnvcXu0hT4z0+7rkVcwdxIexVN6IX2c/cDyyhI
YqWvxNG8ZFA0NgTY7T6jARUZkZlLfrLXW/vhAFpb96+DUI9I5Im8qZVMikqp
GGBS7z3K8xAlCrkDALuC9Gx8zBKw9xEayorB6VEvyPzlKfRdcN/YIzieIgrL
XhTGUoT+G4wZLrQYCG8I6IaNp0PVHcTHcmDxxSy5yFKq+/6beMkH5/LiyExI
Na/dyjQLui15OmRJco3mCsh5FZ1zjtUs8gZx1g3WcqNnSeS66fIznCSviguW
wBl8K60Amrz3jLavU2w003AtQBunxBqM1KmV/tOrMqzKRUpwuGMDHHbwWrp/
EfCZQcRt9rIiBl+xMrCYPBiQ+OPGLN6g6xE3hsADD8+hw5fIg4Lpmqrnl9VK
F5Y+xo4vA7RNyscYL1HBYElTWq7mAkngKLrsrNBva5r6V/6Sm63urpKghYF4
JtTFdRexrgurc5njA3S8F2EBWq6tLbI5m2PVlK7z+LCkwV8EoEArcmqOn4aw
MQmNdAfykLAPS/PJs9qO5NP52J+CFJcqhXeFPnCS4yOTSF6XODmCC6AW4PW4
n2bszAk2ywu7fFAoykXtGKHLk85m6QFpBO7LQ15OtLMCEhYXm2qwvt1xxArd
V5/5JoXvLh/XblZxYcpsyq1xGNdcxaUXYTOuPXbYDr7zaiqgDP3rVtPQ4mye
UqVSQ+LjTotEYynYYzWwuKqOAHyZfoWdB6sl5LviKSNCcvAteTTWa43nMtBI
aBP/sUmC2xFY403YHcwqyswWRZ31IGaH1kRfaEGukoXRNnsMdky+8gV3zc4e
WiYQ9KXC5+E6Pj4Jbd/KOgJ2oqDEqIpss27L7S+DxeYANKb8d2UV0BPtMa17
JVd0aee7zrdls3PM7ULCF4yu9P1RCsmWZ113wuD0bJuXDA9Yp0PDQC2AwyU9
rvKxkczqjtV9F6ix4SQzV2AP+nXgNxFjh7Oxg2TX0AwnsSgso+CaPXv8fJJ6
egLQsD/T58RSDRbqi5WEPsiY6L9XSZE/vRJp7STb431NzW00ZYz5OSk43ayU
VRW38X3lAgsDiFV1A6AsH4OqzXi82Js/t/NffJBCfEsfdz3SPI2xdPT0IbxZ
C2uV670WlimlfSG4WcwTYWXHHtXq1CetYhSgE5Ia664RGHevmeu5Lv+7NWWa
QFuutyaonS85bSdQf+hmz2Y8VsO8a47FvdJUIZTTLt4Zkxnd8G73JOVEDE3o
KCx65g84ni+iWuYMM2CTnI72hB1h2BZXoIu9CEZf6NvVaWnUMmtJM3ZJ35sP
LoH2R40BHNbeaVtst66twTvyM3O4/l3FjP7sfQlfI8PT8bZ0c2A0N/++h/u8
QwqDrLgQRADrzdfUBocvNGTlWsPBXC3HAaqQNnEQpbvnz9LqnPsbxYN1CYtY
H3VFf4ulolWBwONAukbC6RfoQd+DAV3w+NbqgRoYMJx9WO1MWKvcW0rrQZxo
/Uw+JC8seOX5A3SIqD3vBNh+vy8ugGRJr4Z6wABDIFBUksPwkfyblE1NJPS7
LPX6Bl2EMorHVvJl6H3150KL2F6rlOeKkeZjaDVN0Ln9Fgg97rOuYFWhQrh6
Uej6lBTHQk/e1KiTBQXOS/34msVOOLAWEcs92lLVO6kioP1bIRXshaJa3dtT
IvzrJdI3DG5qBmrKfWEpjv5wQarJhUXV93lhqlBxVZWF0VT8+/EAPqrhqNqK
MZdkPLv86pEoGzb79gEcHl+LDn3ub8ZWApve5nwL0g8DQF21YoaxiD8jQaoG
a9i6ooNq/lbBjDVX3xGJpTiFtfTT3NSZoX+/wKLBZaUUSHOjjQN/5p/smhwl
pPCJ9b2tKOTuDJurGFs/hAepouvoMoMfqB3f0XNwInV93AdlUDt6TJAM0bcE
6kAyxMqxz4QrN5wjBNZVtqa8hMI3NrX2LngIETe04PXvQo0qx44vLn9vELA0
nnfhte97YAPfA5SMV6Yx7aFU+BZjuFy9C8ddlZfaU6H9+tQelVyttfdW33jB
2yJnc0nJG4le4L+BWibr2p014Qu9TjAmNvmASjcVNaQ1rcZa7NWcX5ScmiZ3
oFFo7bnznlj2Vehp1CtKhxYrvUQNAuy+RuhWNXPp/xyhs/EkCeovAw63J1gi
bpO6BilT0s1xxgu3U6jqkBVtv2WI2yEVJFLss6tOYXl3lpzxsd/YC6XXFnCN
QDTQD++XXEU6te3aFL1GZ0Tz8CGL9OE47Td5gtoOKgwMGLErQsFisIPLB24C
P7QeBecke6bfeuitM2lVf/rGs6RdL/KurmEjTsPRExPpM2lG+L7HJGKPkmmg
pP2jmUvLBI2rv8KYNvO+jQTCoZwWkZXGMc3/OjBtJxppErHRPbcKWIDoxPoZ
MPuehZPaiOR/UrNdDpx29bttKMFXtIl41UzqW0QfLtNv1DG+DVz9zjtYKumf
5+Zot0xNmFP+mxmXALdghPI5e52LbOvVCtst/TFK2LA9wahCltJVhOMDNpVP
sr0yEEnPLng3kSwmkVsPsPYeHcbcX6UUOIR6jbitJj4V66m8TPVeHPLE/qVp
XsxCLbIg9p6HRu/AUvLH/GGpndQ/0k+Gh6OrlDkVtUZkO8+SD9fJaMMhIkSr
kC1+VmL4nF6fojpkpMD1vLD5VKovOaIF0GK4K7licGfBwNc26xJInutLIXvg
G0E9HBYyWeRWO/ZkWFOmEOICW+jD3vbXjrIz++evZHRs3APCV7BnWHo/yYNv
mzoV6dLsfuK2jg+JpaAcNPWqFmwBN5eTAoTFZyL4RAhuI+IotYSCW+hHEwvH
hnH9uu5Y54kBQ7PwD3B4/GDhabM3UPhp2Y2I50eYXb37zUOQmYd/4NmSXFBC
/GNVurPJbd5p5ZcObHTtIiBnwssIcJWDzoXvR8GQVcIZsUXhyrUv1A3hhcKs
anECYEIFNsL6xayiP0J4cNe6FJgKMyGoO94eX+Ow8XSApTiypGtRd82ptFrj
5nSMLS9vhlH6dU44q92FdjYo0IU8tvBHJXZUO+cTZ4/Z6N2sFemgpOPL77nk
fsWnM1aOA9FG/u3+qHFaxKE5SCzFZ52gohrZvNNvR3NyjSJMT46ubMPsXTpw
Ix/qzKap1R9c2ezWy0t4yf3g9V+sOl+G3m5cUwLOmie30H9/nbFv+gyU3NA6
VbklRmtWlkJNZbtODA9PZIhTu7//Q80lx2YPijKSBAGPb4N+faMRC8RzgThq
rvPbg5b9ZCALg9wLOc/4Gb93FJPTmJEngMIYP7Yngi37b3svqyb8mvf6YtaX
3md2vx2VxRIZ0uZISD4Ru/IYCgkv9kx7mMnZo5PfVO7hkYnnUxyxQPjbZLzH
06f1F1NK2oraUQvXznqAeCE4cy+vO5xvq81eV4xtuYkdNz1H6tBxlOdOQaMo
jiAdT3DddT9D9sTfbas8sovdYOOn2Z5FhB5SxZEWWJC/7mJsF3UGu3q4b+y0
OnuaXrxToWmo4l+GKKdDY3OadwnKxrS6DpieElH60KoZKikejV7FyGc4zpt/
c4AaXs4F5dFmnDHb875NherP3OhtZr5yLYySNxccX07MNp+kip9qxSAQr1c4
/bu1iJ+1BGmnoCb9j1RNbxDVD8VFOD/MC29p7gINO1BG9FIl6sNLslbFdqwj
UXWof0BYLuPLLeTT0Ii161GW/p8h4/3cPtUb/61MG8w2CRnyZCR8sgTyO2xh
sLbeOFr3+DDZskGvD7D8Xt9/f6YTydt1SbtLTLNuv/c1ZyNTq26BsNvUyCxY
En26wiGEgmFiDg+bdfdRePWKDLlmXKPkiGQY5VK+5kDqYgfWxBwgGomBMRY+
xdIVVDjgl5MDOw9Z5iqjsvljePjDeG7yh+aJ/ynM1xsW2CiQu/blKJXeomD0
QaAgnqwqK9QFOe1N4pbtz8w4WVSUJhI9S5HxDKuV57GFd9PCwuhUx7ufQcSw
UqD9ePLV0NZwwVYGdGed5cIPACTprGk3DmD3Nt81B0bGvk0BG8isTOaOXy3l
5Cak2EfeW7VhMdz2TjXCoE8oas7svRtI/HN5WAK2sp6AuLQ7pNeWk9raJdjB
HPmOW6/kkll+DK+4roTx3Dbsd6TkaLEfBeZ0Ky0+7kkRK2neoXr31KOycCeT
uZe6G5kiRU5xtGKEske3VKbeRv0OsNEKN47SAVaqf8HpERN1h/EmmusB2bph
Fx5oAx20P3rTJRZEWBfVARC5Li6ETMKlwHQ3WTJJ6m1Nnk62cDV5lai59Awk
XFVybxjF1JCcMBF2WEN0i8g8oz4mQlSkdb9HFEFWDudQiMEPsg6600Zc8arO
mppWs9g1o0XXPSI2//iEof7VQ8V/aHeeA6tXKf4CmLxQPrp791gUVjREDY6S
uyBk8SQ6VAJCpt65tuOYOIeBOF+sThHDMb+wRj9Alfbd5QmjEw1EIZpDRZ4q
CXJeJo/jDLs59csGwZcg7IAWGwLysUAlk7oKTkLoCxjVFgbbshEn8wRQoNBq
oYP6S3Ak2qNJP6MwykE9zrWuTvaF/RdcnueT8FgUxbGeo9+rZb/JNATIC9eL
uXkCBUPK22NF2nbpQjqfUWXMM6HAmfTSbJ8R5wXrJumdwL6VvUR3+MFhCRyj
iIoeyefVrvV/qUukTQ4c+sqsU1iip4i3Bvp0e6iXC7mhhO5D6302IykCpMD6
8YDN2IlJWWPEsqtCtvRNO/Cj/y9ffJHLIhc7z+yB8wzcEN8Kp8bexs5jCcis
hiEeC3arbHZI3VgQgI2qy80s1XsCTpwKeKxBYUVOHUSWqxI5L+v+/43h5m6A
wUZjghsBjk303CxO1HRKAJ6veARQUdIqXlLsGeipKmn3ZyRnI1v+j3urr7+g
NHBHAFUBlFjlV6EInLevtPithGixRBEMFqLWEAPoeD/+saNUu3fgOymHfnaK
Z45hz7WyNae/1EnkKsAL41dflv+uWW9NFIc572Tf578NyoxuUhurEvWAXwog
dT5Hj7F+k0jJqi+AV+lhK2mNS31G7/CHEdoqhUPOEEsYgUyGlL496HqW3V4E
7KD58v8GKne4qZ09ZtMjSmWMdZnu08Ft9NWgZRNU0AnkK8uQ2JOjPBr47OCN
DX+ZRzjBTV1Jl+3Q0JuKmZWX/9MwN5Ub1jd5aQw/nfur9QTnx2dQrdQtd0Cg
VRnrV0rQONYqXGlvZWZXV7i+nqZkBqMAO92x7YVmUGfkrZBG3SfaBpaJ1na0
h9EFXVapEikMUvI30G6MDSfhVNm4nHg73AtsklERHb8R1v7yWcCEmLIMF/RW
Vfi8zoNTk6Z9uBXVClmjEvjnFn6vmBr1nbEjHleN6XohrNjCHsFUMr88zZMr
pO8Tz0WirsJAjmgrt2cjBhgNCZ0fZn7ZTpDj9I+sLxbzQGxSl6L0h7zxVtsY
W1kcRt+2RCn3UHI1+30do2nsdM00+phLGmMELz0Zafc0meQSSRaHGgVMJkh1
PVuGPX4/wgHleeOnZljLRO1OtAVlZEKenarZKunkKQ9RSJi/iMWR1uz/9axG
U5Dq9Dz4JvrD0b3RpIhbeCqxjIpzyBWc6ybW9/+2s9VjpYe5MbDgHNGf7q0l
aoAmvuaKcjTmLO7GbP5Y8EF5bWFjZqTpmwt7qhrfRQiuySX5GrIvNFwbxN2Y
yNS5Y/G9DAG7Yk2a0FdSMGqpVJo7Ux6WSrwNeDYXbsFqP5aNT8VF+Q16Bydw
l3K3HuQ4C+bS88okCln4TJOcn1v180nTPlMJZEd61oxdkaEImRSSXzsX0FjS
zTkJLs+U8sUpHlLa3dT1wA4hdj7OAGGd6F4s3rJIwECw6vpk9j7PEsDJIZfy
s1PdBzopysRkDYQdEyusZ2gE7n8yj1nRBhAbd50tzCNSO88uOVQLGRbxda3E
+SQCRFI8G/MMT8XQUZDJRVBVTMaQZosi9a+ovDIgeIE9n8EQcoWVvqZoDgMn
lzYllbD55s2aD322vrIx21W26UnIKE/d50FuA4U9hQGfvb9SFsltjl0YDP4V
ENs6YzfNxLOMd3cbg7g0g5sspbmLWmj/qGmL/+oK58icaDY86GzhGywU964d
hmaunswhxkHRYd7ufm7YPPBJJHYluff/+D7ltSmpB+yRctTpYBPAXNsHFIuo
NivzBwBBJ3wDxbnseT2rSWusUBrOHZjXNztgto0v2bjASMg3plcToFmqtgi0
v+VLgM6yK6MUE2ViOCbMkaM6cEqcsju8FDFm3at5d8GyOArSZpOpyINlGM1q
OKXX73BQc+oWpDdV9cYtw1BfghQEVhqC8F00W6FvBKJH6ht+5naAyueK7BWf
dIlRuw9QDOj2q3weMiL++87Y/lyCVK73TPF0WAJ8YVZd+KsUNf6VObkWYufx
xmVXTVM1brQd8iPLVMnj9b4wKoeZkCNXafJv9w5EZmMwAfCN1QtFhU7fndsA
yxvYWgHkMeUwjKMwL7zZjlQhch2bMiQVwSOycCX2ULZVtvHqzw9Y6Q82jtP4
BedSX1RGdzFlATYqvvv+0eiJdL8YUCiEU11KYYGXFLvkPtO3/y5dcp4Ztu0P
VnMxeYzA81siD5mHgBlll6DaP1S30DQVoiM3lawdhyohZ2ALZLsJU0uOvNHE
FUtl8fAmyf+vEjmYTOiRmanDDn4NdMHguEI+bdmaySH1mj97VljJt4GhAfsz
LuGNv8yA9wRUooIgrSgQmQA35MRnFDIruRZG34JBqPMk9Os6Hv7rezfJ/ZR2
UX1Lhcf+HOZX4u1jXQjWUahM6IGNp+5E+Eh9cEYsNic8hW20TXhlAe1eN/Zv
3l/MqC1DP78MX+cws96xfb8jB7VYT3q1cQGM0q6HQmlnjWPyCwI+V9gaZimo
oWNYmUeLjC3glidmmKiu1ePnMErYTYFrX7rNBHCP0igDDb7Fi3RLqswWYJ0V
Tcj4nT2LeULSS9CmHY4DZjVTyWQx1GKVzIa2EMnHECawJ+NJjhzdDjVIWwjA
b/VTKvGunNOEzlRGkGFNZ7bhiYxqdIUFImg3bQoFvrwMsWilIPO00arn3+Sd
fo+8iAsboZicJPHSD73hobTpjTxOutiZn1J/vtWtvEcqhI5KjTaJhE4SDxvI
cEo+MeNyyR36QwjYttgzvcaEihcN4YxwvJ23xaONYO+jDM56HLyvnxpTBXBz
kaCA9tmGJENQKkdbJTTLn3UR3Hu7gmxMhYRMGEDzU0w5bvy4pyCrnT7Eeoz7
Lynuy+c3RyEqscdRC31Rz6rjX2hp3sT9og3M68W9HftBnkFQhOS3izt15LAu
fAAJwv7GEh/QxBz5KbFa8srTq7UbUxKmB/5QZmrhCi7VsIkoz5I3nNK9vJFq
P55FWuvydnK4aPPYhUKwdr6NE2iCiTG9o3zSYkb5aOpClFIzTYpoKWGY4pov
9ii2jQFTioKK24yj2nxfHQLUwXR26plPaszQRWKO8+xNMEjvDHV/8X2W8HpF
r7VWlm3qcHQkUebPv08X5Zr+9cZ7/WGTdO8l87MBthdv4+PNYAYftE4MtyFH
WwRSXpC+6GKPpFMahNrANy7yndMqgoYE9TdHiOXEV0g1jb9226F3SqOSNnbo
fgEbS211LnB2amrzNqUpafNyQBQjcOfbVMHh5kXONlfn4uaJEVZALARiMkad
uDIlF3YBL6N6Gc9VgfnE3PkoMHi0eHaKVPHdaHWR/SAcHH34faLxKMEJkvre
QoIwv+lV/q0zoEyar7ZXunip0lnok4VgQkk6OdmGVtw7/MVRHrtiW6Tq/0rO
Ir//uMggpwg21Wmu/D6XuGVRGKKvT4iJI7bIyX9x073Vfy7V1q6+1Gl5SOPV
mq659p60KadMEpv+lIS+0YAkXlsiIz9wBx93r+w5P+tn8apEdv4loOUKQEAQ
fn5mzqXYdZts5W6lYSBDkBRd6Jhl6Xt17X1LabJJvKpqRXI20fwfSvtLHcpT
Y77qbciC5oq6O6Tv4XjR1z/AYtMVBYFXhmO9rrG0w9omcGQvq0xwSwr5Qe02
gmhRsRlfVhO3dbCoigYchNJY8O8rvPZArLzZq5FNVUvBKMHwtkaVL0aPfXCj
UR3nPJOjZUxoMQOTBpBuhF2u9i5wqT/bTnm08vTL/haeeP+lcFRC/D7XOKtX
k9m0mLyXVgY/ZpnbuwaBulZeFpvyNxjkUR4AzjGPe08/37nRvF8cdm5enWat
xJ+7dNHSPNqg+ndtWXtUXlSMK8gl7uaAkUGvv1RPQALJO7Za69FUmzJBpcUL
QfPYi8mPYwhKrUQ87Yxdymbe+PGyb1FeW5IusEBjvcjquj7h0s/YzzARyAqs
CsESUc3AwVwRYG3qdSgU0BMy/CMoiGIrjur+3aBqLZfukIGIjyARqCQ4lg44
McLxCP9CfnY+lst6Fw+bS8g7VWHnDymlO9SaJe/o66hro3PPEFy/xgANue/G
EHB9Z6YGRiOMm7VwX00M6H9ayREdUGYdLcG7IgsiRY5PFyhbctvcFvg2J70p
7W0xCcYPFv9JASPRcp/hPdUKCmdIUtRZSfK4YKINIrhc8QgbWp4xFpIluYsE
0kxGwRABO7bRHMJBUhksbE9PmP+bL2Tt1nlDHesg+5uh8RBZeO/Wz0+u3k/O
soSX0FvWqqmGBLaWAvgtGvuoa/HDkYVfEY0XjRUPilLx4DOFHSKE1SG03Zy8
WhQtoAKeWjAAJWFzzkkD0go+tfgWiI0hktlF9pKfE7/Hlpt0dER52KeEMX35
7NqvJm/FTZNZBnAkp4VUl9Wa+4aE7oWnMstMJu2VgfMbCsIPpkbS2zjTqKCx
gaEezx/6DewhqV7PIpOR0rSAm/9kAI69Ecdrw2oSPAzyi5KTOJDv03SZLP7j
wm2PmzXueu9VAquajGNkNnq/01ztTSZVkYVp+4W3aOnyTXSrnV9od6+/XPvT
I2ZPEKtspmA3srpT/SHOXsuL3TOaYm/fIyy9kx+ETKeJZT+oJuvAUjPa+nfN
cCPBIcT1mzoWIHJEFNfr7Lsdegjy4yegIh5LaPnBSZHNYX2dW+TPqAJ/BrKL
vna1zKFRGiSIiXkqRbvWTmSt3Wf0umZAUHcliktPF2yYC1jts8wm1jRF3Jko
EnH1XQWMhwCR6Pe4weU+kf+Tg/A3V1l+VXO7qViueWwKtkmtWrsT9wgsh2qx
LQrGk4xX3Gzr9V4VokCWySjUfelDorYGUngqpUP59x8Z0/817WhCJvAPIBCQ
2Q3kzmjODvI1ddjM/Clh+1/vtwb/ACGlEDqCX9i/sfW0YWE0nLwWeeE2ehUN
4h3uCkcRJTTiVy24W9SoLQ6TpLXo13ubHXJ5/je8uvDrwXk4dOFPRD24UexX
lQkta4tiEOVjfJIfCWD9UAaa4Toee/DyrSgj2yjrLXjynTTmUvlYdobj9XVO
h7VJtdPE03yJGvNxFkdRrbJKZPHtFUhxTJNjWUbfvG4bGYLxRRxzV1fy5qij
3eLIIoQIUZDXG3HUI6CiAIlmsFqdqnn52vzHaAZdoS9S1b6o0OTgay7eSiOe
kbAU9/fnuj66OPdS+ktTRoyHbCRF2IoTUJN9GArXl/ts1XF+8fRhOu8Vso3X
QC1yNzK5U0sCDhn4M0WG4y+hskKIJBGWXpK1855FvwbDkWLGETNby3wmLGlr
xIsgkj8l9/1eukmS6pWT5/C2vyBlaAYZJTjPJIvvveI4tD5z9fUAlbDsWEPx
9GMQ7ESL/Xw4CR9pYu9re5EECqmHxoHSYqvV7bwsh00JNNGvFKtLnimIPTya
td0r9xJJij9pCTuh7tb2wxI0GTeR95v7QLe15vBJHQxgLeMjDIqvvEIZbNSu
iJuiIfBh7O3VQZXHnEpU5h6IKHgSBqJAoJjtRxCAqr7btBWERXlehnrGtve4
/M/1H7o50miuy4J23BXIJ3cQlRyjfiS6sy80pD9C1lB8tGfJmJNmZefCOMA4
pOjQw6ngLGNoSaj1lW/4FQla6eooezT612D6SciamB3coI/kg4pSd90Z0UmY
mimM3or7fhBk8rQ/IIKhPeKkjtnl2qC1f9wgITvZ2/UeWHoXmgHtd2PJkKZq
Pf22hBrMWt12RWrXi6qOCUN/SMrcebe+HPlSQhzX4TJ6wUkU6jJLwcdaIToo
obqym4n0clbWTP2SqIjoWsN7aYhdVn01jqWkes5Sc5CdYY9ZBVWIHe3ua/1t
OkjZybGQpJnN6RRdqD5Qyh3eHrUaQKlx0IGSjciDJqcVjDXRBhhxlzXTxqmC
6f1/hWIk5ut16hs99CYCTBHJIPjDfmoUCUNiYO0c8Mo1X/ZI5sKXYMTE1uwn
WPmU22fzUsCrwfMxJ4/0J5GPkQlge+hBFwWefVP470TLATt8sXCPUE/AaTry
queCW8SUCqUu3KwQExGuN4spleZKhX4Pa+olLXTBrw2wk15flibvPL2oScxp
numoE3NPOgFa2Jh6a0NBLIKzUBN975J3FB9UJNdyjpM+ICanrsqe06u63w9h
grgL4OGmg2PqdLOz7WQ/3zqQFfztX2MT0d8orUZQ0enITVLbn66pef7UvaqG
OMQiEGzytskHqxYFCutR1TdyQFGMKfkjBcjmxClsg8zg/P0DBEdJVNWBghJb
mx2USuxogRPio8CGyaB3MF/BZ7JENEr2SfIzLQDUdXhnF4HZPwM9VV+D9tFv
0QebhX+BQgeJb+ZuGmFZxeXPjnBGKhQ7kgiBr6SEiwcYEB/8spqoL6x0uDsu
knP69QVWAcCUHcn0C4etbDoKQZucjRWg7vy6nDU21G1zmbKHekAAD/0c7mZS
w0D8mFuUjPjFJDGEltdcJXCSyUWrglOpmk4Q/v0MCtS4N288f9kzfOu/xEtR
waLc7EhfkzVpzFkEe9lfo2U3QjAIONBAFC0vXzp3OEBDnl+lqANTTgep91VR
KF8v6po6HGqfUTKyHSiN4MX8BxbSXVY71MNWKTSMIY1RtWTfJTyaQG1OF5NQ
pvOFCMq4NReeGAUjiBIgouXzeUJmonhTooOLQqENJPPnADfNf0Nss2hJsjm9
lzQk6jdrr4P/NgslXq9QaFCMAbzSi4hDwn5H2GpCCla4RXpekdepUwjgJG60
yuHrL5z2yDdpexRCQPAU85cGLskPMTUSIdy/ge4bvMFFUmvdnHvTTL5eWePS
PZEkmhi8Hqh79SxDyHgczmGCSjZbyQzhCptWjzlmm4cTXz4HfSbN0JpVwbPF
GpsFlVtrpdFb5GtO2heEFD1YcuXwY2QomjgT+EWWIIr6VUk0BtpcSgRopr+a
AMk4PjbALHZ1KjyeM6YFVwgKhGOJiQGqK/qLm5yAyPwWQapWtKXvSPI0R0/2
34qwSoIPvUZbh801MxB2SEvmmXut36ILH3P3hOG12mDNlhRqIddz7DhBbMNh
2WE+f7GeRSfrqMUVDrGYMuOkvzxPX8TTa8tJLbIZUj6Mn0XjWOgy0Fxsyt+G
LEAO/XCNHtzwYlGv+bzOHSQ9xtZm8tz1mglDrJoiL30vmOHKVAWXQynQ6XCQ
WXiNpaC/XEPPn8HqFwfPC+J6mFFlP+ZYTlCjnm4o5Q6kxnfbWTQ5HcEiG5Hz
orAY3rVlt0uZMBECoDjtgzcUd0EsZQT3abXVah4mbgeMBjkbg2LEqbwZE4Cc
3DIc4zF43be8P5xXSdFoM+GIEbuaY/9GnhHUeC1vDd2HxLy39u+mgnUZv/wh
8O5rjrnBgd1Kzz13//jER3aShRP82EQKtD+QODynfoW7vFtlWNpNw02JsYJq
0ODmgitrGM6LSPkdU7qi66PSa2vNUfkDimK758uu/RynjpnUlsBgRTHbD7C3
rbUn40F9u1VCeKxy1GjrxZef0odpa2Mb3qA0wplwYrSEjxaY1nkm4zioWrJV
AVTG79lwcOvsPCqYA7/nXSVn8h/kQPbj9nMJdraiMYPRI/X8oonjVB7is2TG
SPyJUnogYqrpPSmSdgrFBmavklb83X+VR+ZSUQp6Y2fNd1N5bGmogB8Fwo48
CIt/YIG9VIqMJiq4R7DLSjgmZs8vAhYc7U1/Ii16dGMCWCAxcepWNOebqWLh
QWCNu+nUpHSGqK6CS943on+ZW+vtVq0e5OWGlsOwxk5XuOfb8jnaWLMseulQ
ThWv8Nk2unDqhO39NwbukofkoMuYjfyDb968fgMAIQV6YLZMLsgKyAHQYwNT
AoUkXlggAba7ltQFAds2agHTe4EoVmuIXROihzeaT5ub0jLyhwa1ZvxzzgPu
nXlqQxG4iGlUGXrkJypwVQihMjDhgVBSUTDS3bH/2jcqLo+YuNS2jwEKu/kq
MADPFQFvle+6RULOG13XZgDRKtZFG0wUw9hNgIb8xZGy7OOp+WfIGfw6fo+r
yoBt7M83IhQH8wEIlc/5miL7sSJ8F48ORxus/k9TQfExFw31f+qtFbTvpuWc
uNEjm9ECf4KoyPlsUbXYuBZ9QlpHBYkW8cYd5eMB3jjkENu3X50gB/mpTfRX
HE7zyvy+Zq9mnI1Phplx55AR4Fo1Ud8ACwsNofmHwDsMetuF7s6k40RVfZUZ
9Wj1pA7gDnkkLKAbTcg034J3eXYI/9UJNvQdPlDEg7BOEDe1bgB70jLl2I3q
gpKMpjRnOOWjEOY24Ex1XiOvBSPyl2qhtcUB/xbq7qjJJ/TuL04+hTZfCwSh
+m8A8DOWwLnhAhqUGBtnv84O6mrWSDja0P93P52M2hR99kY4wmh5kGYnJUZo
CpIAtXITVRz8HkNcwU6do5qrKEQb7tgj71Cd/XSxyPcerZlYK5iAa8CBPLH/
pek59VGPRRV0uYs7GTtxaJXWNFT7o3SCRycLkGmMcuezq6QbOp8Hb+gVxADo
wBT++x2O0Sh+HpXj3oOHOk0i8WR6ej5k0jYFKIK8FWE0zBEKpHXklPmwBfyC
CCNO1tP+x0GUJ5csH/JPwSA3dDo2MMA50N4IMhfrrMbIgX/aW8CEGj502s4+
DqvDC7O7O3MDqaVVQZ7zOkMmu/gtWElJa4WCwtFPBkL3lM8Di3KUDrXXfh/f
SjAFItV5N012YdBf24dTf0JgnjRatY0K//S86R513kCp7AvLCQWQf4sjmY3M
tnmxjJ8L3K63L8mIbMpSF9ke1D4rJr2YNIAreO+lfCN/FTqiaFTwN2XWDLfw
2MbKDecrGRiPhAjPinAsnRUfmPsrRuqaRn0n8HWbpzcympMtiqtcgB5SOC2v
t1eVUhrn5Qsn4x1VOSiQr0vRqSzYRc/PprPSKHS4j5Pwem/j2BMPjw1/lR3A
W6EarxtGxPBU5l0+1Bi/1+v0h9Opx+RgsKm0FT0jyluzZ9g0K0WR5mnv60Rl
2cwzAZ20Ox/KIKf8TnT72TwI8zR9jS4fMoegOcjG9PdPhdXv9hc7IZjL4eQl
jHKO3XYvqTC8AB7sMMdYXoW45g4b2P1gKlZw+p2i3RFc499Q0328LQrN4Qwp
w3UbMdm4cqWQpeTYiB/ciM0fnuSAkqrl1cV4fFlY/Ratcx4t0w+gOmJGtYAw
lV2c5YX3xA+8Oz+Yhd5dfW4wCNahhOi4UgDFwpQ/9Ef6uOJwRO9hFOKwiqom
6SHP8Ngu8L5MVxGDJ/mEyu2SXpyC8gwzsJfW/ahAX6MzVm3g5DSzFjpyvbH9
205LxDtmEPFnMurbDP4dZJWJ4X6FNbXpdh5+w/Gj7G6GEFvru1/V3RuUt/sM
gaSEdMKMk9bTxb15CW3gTEy/7LJwwGvP4YYntbcjW09Qk0Am12lJPQiDzzu6
9CGdVYz9fwOGzd7w06uWdLe/4UzMvLAF6RHSTD923+PbvEUvU2J32/2AZW4M
WtBFo2VwQUW5FM3goyvX/NfDIw2860fT60c6jfsgkv2ywN/9aK3EH9eZFslo
7YF8Ak2SRfyg1vqApzj26/3cvG1t2OJE8WuvtEwANUpeEzNs1V/qNTVGZgu1
sTPQ7XvkZdVYTI1RRiffDI3t0XZnTp/+nR6+66tLETWqUgStVFFpJF/9GQIK
yB4YaXvyZflbNS3mwxEoiLlY/LdWf1WK+6MxCBweWJmZE7z34eeJB9fs1T2d
snxtDf30rpChYRP3VRetEatItkCLUV4+j2i/cbYwNfAIKXR/M6TfG0s1vreQ
nUHFCLJNwUN+8/Ca7saGsUfSL23lr+tkp8FyR8m3ykxx2WMuh2KOfekhPKsI
Ybq9z7TRuLiNvJP8V2uMovg59ofq3q8DYnKgyrd8mY/PK7Fs5m+t44tsAWat
nCg3SE5SqVCpZcBW6YHQrV51jTYNbYr16nykcpi7Cj525l0Py0bfSU14liTm
y7efWDZOw69flF59elSHy42TfaRcJztkWYNfeujLVQT690bTeDoAgQXyckak
k4aX3sCCx1z8ZMC++CG3DM/TNgW1+jryK5PWww/8O2FFfvGgSOUatY0frv/X
Za7fQHLUd6tzRS+a+2BlI4XVeoUOIy68BUY/aNwBOSJ6FJ+unEJGNlu8RqwP
VA8PGPXXYiZcd2klDdyc8f8LGlhbH+VUA6YMZi+G57O3Y4np9ydHfy6WGtUT
ZVj5sXAXYeSiR+7Zae+F5JicY4hwM0vxUSwLlYhOqxKnh15kWuA7q9N0GYnL
W1D6Kr5reihj92TUX+PeqnkI2TDrAABghW5qt/jH3QM7ZRx9eVC2PtU3flUV
NgYp5uqnozSjNWHqmYwg1kguAFj3hY12k7Fxi6CR10jFVrB7u/RAojHcPWwp
LyPthxplyHfbIZevFzDv/gc7TC9Hgwqxdic1JvA2OWc7iFBJwJDNudYL/eli
jdMxHF2ACP4+Ws3FUT2+tMFOIHwuagrZR63+LdEiMRwgJhdb4iu19AHffG25
aMaTaclLFU1tr66KZgQ8r6bK13FnR8G6kVsaHBBBARW0AesXbX+WgxHVvAFq
cs7PJFMt8wTGB0LUZBTvzDfkWrKjw2vA6mSDk08+hz3HcpVpHiwQeyc0H+EG
4PlbpWvPHK2n2OJWgVeu2lOb9eXAWrEWKq20XGjBlI6ODcxwAaMlcxEPYiIT
pybjid27EqnYEvo+lHVCxRvCuC/4+xnw9To9TeuHCu+CRU452ORnOp3guvVH
T1hXygYPymrpXRD66ZLfe650t36v+WgHi0haU0uXRzTBxFPKGqWKiy89yEVd
NsKtKvsGdE0jL6gjOho47W/07Gw1aN6puMpF3gRJAWcYgOvbkPCUFmOFL2AW
ACaepjkAF9Z26apAbYIUITorX3dK8lZYtN9lEHZu2KEJBGo2Hoal+vZDljbN
aoIW+Z7o7R9vGpvfQ/DidAmwPYuapXdVdj6RYBfNRbn9fZPRPriYruzbSgHN
GFB13ZzGdgupvPON9XO5o2DHKtF7JpQtOiViUkhWITdwENd4wz2i0qIsviU/
qBOytYNCL0/I6/SuOL0Axy4IufyduIIagEWG30ETxvwx3eKKSuboft+N06FT
xKY2UhwpTMjPTzJpzc4vX+VhYD68SN9A3nD136L7G2TwVCO4nvCmvNs5hhQF
aLsYoxVrk63pdtm6/SYlzJfl5CThXc4KKYrse1w2sFoKmlVz8Ldex88df3qC
LnP0M2MO9hHYwESP6R/cd2HlgBO1wLx5N0MgZip2n+II78Mnby2WZPMHX3JT
8CIQW0l2FM6HdQigxdrXuNl282/QWOrQQzzoTxDhkG2Q8T2FmlOwaTs3aO1k
6LAzAQHD8PYJiB/uEjSyfgUhHPoVZfDu/wUzO0AI5IWLXYZ3Nvopf6ZKcdh9
RsxqQfRA7vhnhc8/yU0GIN9FDN9OQx3MFYtBYVobdl2i0sL3E0avAyrqR2Gh
jb6KMh2rAXBrt/2PKstynhzfIFgXwCpFv6jYfc/jhzHFOQAqfbJP/NpsOTKV
KpYh3DivtR1O7hA7klKaH7+NgwtKBT10BH0gy8/7OdfmEM3qhPkbHmq5QUna
8gcPLSkdUfMeGU4N/kxHnBOJVQc8/PodPWb95ZtfougbACbvlx2WjOPIixtB
RsbMyKnxOnGyWH/L9PQk2Kegs7ouoRUcAc7rkBBUsyORknPnwHm5mvFGpUuS
IpFXnOG6Ks4567UsKGDysXYhsbDJ70EBlDdpHkQiL7ix2A5ZY6PGCy0uuIPx
Jt6OIJveG7u4WOsKAOkjQVf5jxIQL+/6OGPrM7xDCFjAJHPtoHWGrLnvSL2j
+0om1dsHto6AJN/2rI3xm2tldDogLa/k6oamX5j37ZnlzDtREYucSAFmeyuZ
zBw8hu6rbuoDNlw0DdYnyP+ztnxRq7XDIflaMxxLZvfVz65TcDY0LJa0TNek
CsyDbckJ4sRd2duHkljb3MXsDfvepNfWdaczZn7fHeGJFXelBa6gOHmOtZ2B
oWS6FdqDdQ9vbhRupREFBQ8zsrkYE+uKlPO9qNqnwfs1gNDp3PUxpIwvjkQS
tfh0X1taVHaldlU/kleIMWJRg+VQNQoG4vMlj2eq4V/BYSYLJscO0f1uOd9q
FN5nYFkP9PVtdcaMYWGyIMy1ZzLHWgi84vLlBQ2oN4DHVHW5g2TISB0G9h2R
qxbTXOqBttEZvR0PNIl86xl/UnDVDqu2TGn3h6p/qiCHpf8hXuTAWmWpBF0i
J5ttW6Ri3MAYUsBbvFiPNgO+YuBwpJiuq3XSA5Kk8L4Cw6EB7KcVgPvBQ/Qg
XwQW3SRqtm8R4jnsP+EcmmTKZ502bMWj/pm2V88K8Zp4y5Mm+iMTZFvAt+Vg
eFY707IOP67OqkEof/sTPlyJfmnWufsI8SnIJzjz2vypqc6w97/dwAUiLLYa
DMSDCMJgztJOZGBHT3Yl9GxRH21IRxNZvzJ/m+TnpSxWjJn5g/8EfZW4l6e4
I+zOhwj4Wmu1nLb6HVacy63PQaQyWbMg0V8iq7ObyWbEkC7YPkJcDuuJJp4E
+5woF9W6vP6mZ08J574RlqhTtkWJhy5LYV16QKJ2vr5GNy0EjeDGAOBNlRnU
5puJzeHVgm3D1ZOTg/k2ZW9fnSRSKZbNJEPptLd1l8l8ju4zlsSPTuLMSRpW
V0P9K0VqgezN+VmIBxLZt+gXX++IQOTXsqd2pOWmeeD9/kTM5J4EVEsRlb5F
6/5NkWtuVSIu+IPOUK7C2yyMvnClfljtUz/+xd+X2c7NCqQy3GiGqQMds7tJ
GdK9RERZHT6/95q+plthtswhRLjdiVyMvCHLQcM+HPKVB8wBKlrp0+BDfik1
QI7wbfL7ufqlueDubExMvbRMy69R7v2vKlxwzvVjqI3C22fkLrnrgBg7SFlK
+9kda6jIGuljLq48QZa870f/XNrM6TAllwprJ+5vHIKW9uhSfaj/Jkd92O2i
8sI7gIFxEYWjadSjn4FnXFzgl+xkNeTOd6Fe5kCq1gkbbNuB5FP0JE8rWfcn
AFyPwptHSB6PcYokESGSIQWT/r1esdliDMGsENfYIuFfSNHqXlee0lZ1qOiZ
KbrdDY5wpOMNLEXB4QJeJcMLi6tbNA6FtGym/BcYEKVW6NCkmQs/0SjSfET+
1641ykqi0RrjryI+rL+LhLynvaH554BOZvMHkK2A6R4ysnCuiHAXH8oIeupn
YDYPCg4+9ONiPlJsVyW41Y4FOCZimCe3F0gcgIyEOyb+gbFBj1EzXwKFi+O5
00ICtUnMaNeq73J4XZJC7ACsSTPhAONFgwS5IUnpZ9NlqeLhCcWbp31psoeB
fAAejtZLrl5YalJ6T0KWhT8onrgj4pR6uuZnQ109rRwpuznAyBA9sMJ73aga
mUWUMg2iszMcK+YODI08Jgv+yledg6Nc0CHZBnPFaq/FzTjAJpyWhpe/3LBX
eyPzR9fC3B19rrLKy+mKKz2IhxosIEoju++3f2niS5S1hkCFmDUJ1lFicOjQ
lmsawXFw8uDbiloBaCdICh9D0qCWoFT64XnIxDJrcXRcHF6ISMI4o53ubnOW
SfcuK1aE18MigJOd3wNMLMm7hnhZ139FobS+kzubilgaX0as86ROZZqEr+J9
GA+Z/s05UInBBBMKQ5rAwwnKQ7DMhKMAlVERJPKZTlbokwraUOvbQ6g5RylI
TeipAwEOQB+Wwga/j0TN2wbh8JOEW7zNYZIJAQr1SYP6xUmWhXmRuUtR8vP7
1wX/28vg9l3Fi5E9o3j8g8+3Is9fc6SGakQfPjlSYPyp4L3dFzkj+q27aoSN
D+XDOGykCG4V2oBBEtSsfWUAZW/4/8sHu8H/7fD7Q7UgDgSeX6DaakpnA/JW
g3clWxXvrNd1/OVOLLYKM9nqJwD/4Wg8FqKzBe864ZkNLDmgUdbKeazFe/AF
B0+TYzPxqnAkAFzjKQITw5zhTUHo9zpplXETVfeDAJ/MmheQDmUhqisW3AgS
m0uOeFomOKGeGONynDLJI4tfD0+9QfQoK9FYXfnz3x4hyUdqpFn/q56ke4XF
UQIh33+myxCp7/k/iPDNybZGwv5fB+NTHUIgMUwsAYIo72JzULemNN9w+ngt
tOiqtvSsYC62lugBvFx2/hIoUxx4yCZ6XTR/zvTPHvKD4IvdkR2oME8ZWfMN
KB6P92hpo1ViYL75esyGi1JfMbctuC26Q4kveKkHwew1fnPewNhvDW5BmI38
AopE3lkxRJ2rfwlj3h2vjnP2+CW9OKNfJvFCvafUkMja4FfINYag03FsdWqt
C4k28HLFTbDKzCyP8PCgMvKP2eYQIvYhfJMzTM7/HUAlb2YkfBTY5Mrxtw6e
A1zwIKBik7gPXTvJstN7qcXzV7Hhy0lrqJmcVFUPQPumZBn265q/TGGXGJTv
TiMVq/ohBkEgkQcD2MOJECbrDvI6j/bfGlYuSl0x31hPav4///f0w58Z2BWM
9/03iU1fo3Uw7t+qD3XAMbMxCO8JCH0bWEBuRyKXJJ7Zx8nZkvEDw6QFgd8i
wBTGL8rI17JOr6jTWa6TPTl6fuohltlUcNliBQ1Gz1NNh93QlRxPuLxe8fbA
lTri3gtOfRCCc25iHmj0Oi80LCGOj79AsAZWR9jphQgRSO1noAcEpkyYEWb8
7yZguXC7gXv01Tch3ls0EnQgRdr0uDUhLh5rZcfXWVyhiBpbI/+lT1KyISKC
U63GypIIGqyTck0d7GKSx7iWahG5H8gJkalp4kAE4Sv3Mxt9KoZz7bZAVE6c
JDwA8SYVOQNPp+L8stM4SndQ8dQXU5uqFv+fFsp6CqRF4u5U8EvYZdnGd+Ay
Mxtbem8c3kzUD1LYkVLP+GPwwuNXBbXrw3kkjQrdWGX5JV91h6GRp4xjOGUQ
rEYjTlt1NYlV0rNwumaFcRXNPCJ+dzepStolai3FIU+4z1yY+FMz6bR8qgts
tqNqG3+rQeUk7nXi+oDtn195qws69tLn4fktmcw294FdKATKDRje1VxH/GDQ
gOmcVdWSwW6qAl5oL2gGtptrX0WMyLzJwER1Vs+EuGkkj07Ei8JqFbgm0Uh3
/Wh0MGnsi6mfZ09aQ/ksj1mTxp3KsU21kkgVLO51MxzEsSznZMQ2wPAxtRgD
1eNdb9EOxzd92zAAyRjUuhe7+BbCWAf0WMCOvFUzBovtTyxldb9zP5dEGZDj
pnoYxvFaLtqKutn95K4p9O5zB+Ad3KLOno8PFqCO7HrRz+uUtc1mYMezdhkS
1bjOKCCB4Onxq/BW33op/WybS5dk+b9GYxUz/FgezAexp05EPVZWQP0Gurtz
uRnCs/RK7W6P1frWEm74YOQDLs2fzy0mtUwhfSP8HCyVnPYK0FIjVqvLlM9S
if/CiyYgGnpSSjBoqsFnvHzvjJZoTVXuv7PQCINVQiBcB9jNxOfEnQRCh1Ij
HFiHS20Cj0c4+n2FDZBFj4OrPfAcqtP4WIXklrtFjl5olmmBKzAYu73TzQou
FjFw2bgmdH5mV1mRglSPlsTlFt/6HXs0Q0Mx8VEhDiEsOHZZZqJGZQh3XmH/
qdh8nR5aVA7YdeKuvDfxAuGOOtyBEM/MRx6+qg74fOUTt1SZ0v8xr2cgrbck
guqCzuJPZFW84zZH2/BEzNEktsgrcBF+HGNyr+9TGSiCIOhUf7gHQpnTtPCV
bOY4gLYSORmnRkc5Bhpik5ZSpoasucQtJi9ke0uBLWoqYBJSl31IaKDSSngF
iY1GbahXx68bg+TcNEKQgZZUZCjt/5srTvT3kEWQe856UjO8M9HZ7PI7RoDm
XuIYRNR7oVYP1FbShE9zB15HywPbMAF2o+bfEbRVc0XnMKqi6kzY3K66wpnO
w2FDU2HWMHyGp5Mt24Ph4zmlk/Zne61MuNSaZl5QIlKARP+mHHTPofvIHVk8
1Eh0WqBny1bJjSw8VgZIu9Zr9HnOq0NowHL+wbp9LCY/kCjjXlwAQdXM7m05
h11g/7SQO3tm7se8ZhwwEQ5QZwnOXSWDcbEFJSkiFC0OUepGn1/jiAgZNX13
RjKgSjAIX9CrHOHVw91gruIjzqHJ6w+YGaEPLJ9FVHZKsR91JPfqwBcTBbAN
bOKTz575iZG3k/R1l8iIofWTFBdFaRpkSTrkDtNrHjHucjEDwR/o36sph49M
D753crksfJF0/6wzXi5CKwyu67Zs7EjIattKPWdSzZU6XIOwsrbJdmeS2kHu
tOOXHhQTcXLZe4wBxxyHfIXvhbiC7jqgTSW/P768OZzahLnzco6nal10bS+H
p3wdK8tm7VusxOsyeOHUiS5VAr3ITY1DbLBaZj5SKG6UaYCANqIvJMKIEJxQ
adH/XnF+9fa1kuq1x/XRNpxMGLPDAdNscoBeoRtcP/l84FjLOLPMCTrB8IKe
LlIMw75XWnC4ouePZW4tjd2NFTpQQeeGFAwSWcDPKakRyPXNqmSvbTbtFgzk
yklYQgdQ54XdmyacfjS3mbXBtxdZFIobCP9BxiMPiNvS3v3h7u8Dy5CZLXFY
4M/joLTGOSNsJiD821M86gDN2yxfSB3lqBfFg/3bZVqa4JrxabNnXoz7FCod
sX01hzpMsAGRr16AWHHr5XnkbKvAoJhxdsqyhYQiPMI2uRXfh9+9o3oJvY0L
VpstYvDUel23NPXmKzlIApnAtmchDnbiILYysNwGQhrKq4xgG4R8njLZk2MH
Bg0jX46ClhfEIKKjfnW8OK6VNdJrtpei17tZflIKnlA+D8ZxalcGmMvVu+V+
53eJtcSa3VxFwCn1AUaUd6dtD90fFHVdXgXG/6be8lqgLeJLkLIDTDRH8d5R
oVXB6EiwumX9jOB9t70m6M4Yf9lVkdzUk2fbpK6YG4dl6VVCBtBsL9mLVlL2
XZn0UWsPaocNYuDz1nKK7NnjMPcNRy7GiRGdmHTGECFknK0iyVIWHICTdi3R
eZv12hLjAZZI68W/I239HfN301kEYKnGJcrgaU9IJ6r4c/3GzZeo1Xj8L41Z
oVEsbmBt2c3oOACSMAKJxphTvhu9SW5nfU62VK7DwewrcoVtkF/TgxsY1EUP
HjXXHsF492yOcjTbl4Hm58pQZjySPIWxtLAQYqIe/3fr0FXtzurMarUP48uy
JLF46v0pF+Ct0mwyJEUcVFEYUed0YMJpH/lyu6nPWxhjUUtwVKDu5IH1bQaJ
fXVtXbXllIaGF43sORHEeQmh5IbhVy/XQ/fND1eTnd5si8Dt+LSZWsJjwTC9
metgimgGHZBFY8ioxSTgmWf58nZd7jx0d06dZrgKWdUYWtfOmDudfqqmSYVx
mcjBb6N3Qf9z7AEdUmFr+kyI/jrkljvO9yP9v6qy0EEkV2yorxNCYbyvZHPv
n0V5R1MPqebfEov7SZie9vgYr7e3aMmjwXpNWPS280z+K+T9CASXysTK0PHW
D/PSwzIUtgNZQm47LVdUPPsOFdvTG9pCeWk7NKf3qH7wBFOD8s3EYjhqd/HS
HFt55L4RoP9Z98HcvxAUZoLCkF/dAXhOxaGbvkODJFpt7z1sNuhUgyg+P6mr
93ru2+CAScPV681b8uN6UHhpeBUa+/pIhEXQ+/kfGuaN4dGdbMkRMTNgdOSz
DU+uQWObli5Gx9/qXGe3bjgCffuaxi2pJnVVSTcAKRmC1Q0J3T9RmeONuDCT
Q7ENAsuiORGgu+TS3ujnBjr1DlE+wQUbZCbEv1P3gHy8OvHQHBE7bavB0boB
a0S7BK5zhJzt2QRnIxdKVWm+cfrJojVmhxnALchLdGDjqFNfCIYGaf1PsO8o
VR7Ssjtl6LDwRbqSDbqFZpX3vnZPfDzFJkYKo7WSmXPUUZ3orjgdp/daYFCi
3ajX1vVdXnQGIc8E6Aao+ws0HW5LCq7/pOxKzSpIjb1oMs5QSPw8C9twH2Dj
0xSg0tBttSs1exbKIwS3YGR3Wv5dKBcZYHNxuU/mtAMqeP5WbYptS1ihOYeb
0t0JW8QP8Dbw5UAVd7pLCHA1UBbrEIPaOLuWSa8JiNl96BVVvTlfRWer3S8L
zpKMXlJ1KJzx/HtzMYM06yf//QlYz9A3wuxsrR2rpcsN/4HJiSE+a59H47dc
q0b/NJsTKoqkkUyttDbGEaWb0C1uo/HQaZq/egOZMHCdMAoBaVX0aY1765q8
Og72sdxHg/+ytTAgeyAT4zNKEzo9xLqyv9Gtg+hGbCIFDknm7MPkCAuYr711
hRy+xuM6S+PRAp+2YK0wxA5IuPWI0UGPMysJC7ux9d+s0ERPzJ2BzbFOXpPJ
s9bubsvkP6VTgCqtIcSAgJHCtQl5YrJbHNyOEF4cTJdWocWNe5ACarBWZ+9i
IsqeTN9QOPB4bW+UXWLjVOyRfd+gEahEJZFzd9NeSqrS+kRmrSumNJZgeIGP
t5AKrW7WLGbWseT3pqhGhUl+effRBEwo0EJ+iX8YK1Bd6K/G6CiQYmOdHhSA
pfpyJ0zaYHOqFjHQivs5VGCmpzYWxP6FgI0oriQaQOwg6HQOwS7GTWhiO/lE
lwdja+UbCIzldq8pZeOdrO/7L1h3pu4=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "cZl3+z0J02TVIcH2La0evC8ZU8jd4Tuna8DsuwukiXDpscNI1u60Qb+Bc10ZOZqqtZ4tU/vmhVv+F9Ysjn63+ggxQTfKs2i+Kg923+dlDx5ogYUMnCsiUjNQFT2K681kKnmkEcWzfeDuIZUQfL3te9+bwCurNMuLZIKNyzpeL6wfIikv5UkJ883l6EkRUqZ6PRXqY8A29Rf0Y0sxDVqm7tAncOf6le4GAj9AGwyD1tov5jIXPKz2exQK4suoYb96hQB5Wn+tOutLW8gSenNli6ChbWPeoJWG1WYFWL1/e/gFsknUO69I2ifXHoL1WVsfbIej8bLWwaD7qtZ8fzIV+kdSUKF94SneKCJKu3v1UfXkpylYBeUzhaoZVGzKaxYqqxXVoecwaLPxzOcQUHDMG74N1VHHkww7SjhUSuMlPjtOkGhXK6jepQ6HaRbatdVaGb9zHyKHXYgBOmhlOaVUQDFYkY3+BBwngiT3EX+FMCnWcE/mr0mqjYmHHcpuowY/EbhqafAIdZpQPCi6JS/ggTu49bliPWklltxjxlcVbtdAai9qeCWUnAUBLxvR5bpaPa2NCH62jf6UCnUGTlQkRe55SwjIeWshYEVEiKZ4fDRoWmLK27Lqg300OZIg7nICADUQ+ozxwtW53Wbyu7Nbb2Vmg5slxnCsqpYZB1iSxS5K1SnRvtpn1bY19k7+FP/BqXTwp14ZUbV5hrBR7zd4LWRLx73c7V9SogXDW29rx9R+kK/NSN0/SjkMUU0dj2gygl6wb0sIAPyjBxDOzC4vbb6THtIJvROch5MqrCNCIlP0KBxBde2yb24f1LlN/nZl3F7gYnyK4vPekJZF8EBVsBltn0wUB+Fghdfwh2/1aCeE80jxDccL+zQFqM83LeAHEr3TKgoFuGPL3V1IAQPuwD70BS4+QXekR7l9nvUb+ISlHYE3o+yKp9QZuWviODJEFR433+ITOMvoCeHlrf1WWZB0YQWXYsqmDuo0f+IBp0d7uHFAkM+fGMdFDDDDvyRl"
`endif