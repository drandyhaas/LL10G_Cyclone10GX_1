// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TKoT6ku65xV9FWZLeUejD86lZlfacW54ZDxaOxhgThcgoi5nvuN71eeyyzmT
ETIdv1hD9xgLiM4v/oR90hyDQzpNyGGyjqCEnROs7Qgla+VlH/krfjHeJi+c
NUKay6rM0oj/AspKLADwNq1CcDWbCJPhbIbIY61Z01DjpGy6nJIjmIlUNW+8
+S+pViSKRz5wTEw9qNOPVfa0d6VZeMfySLlB19uzyVF0jwoVmAQhWh0x5yqf
KyQD67+My9+qwz3i2jD4fKuEhOimwC5ftDbByBfdzErRluiy6Awu1Fk80D15
aIttSjXsCmn+/PPJ5a1RSowN/fWiUzkeIpf7wVo/sg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZzdJ9HTvHnDoBSGr0rIV4CMcysXLiO4n7RDbSG9GLfZupAVRbgfowUtYZ2y2
EM0Li1znPA5Gl4AyNnxv7IlFAfMxoHmUDlH1gsBfvh+T2MRM+XFwitT5LHOg
GjBAq42jlokpDgRd4gQTKZm4XwHq75I+LllUNm4nRaIgnffb+fnmOP6ZPhpn
hYPFsPItcci15hUrEhODfzfudiQmd7zGbVo2jRgorqx4CQw9yhl3lHYp75aP
KakrTy2YrSR549OI2YTjIUBEtj+e+GI5QDQEMTk4Gh0tvEPxO7b1T3ptVI/X
6qAw5VBBRxqO9f24PvialNiqjHghm72Aasp24CpU8w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p+sO4WhAcybKhpfYEDTmed5Jh4IvtZZh0nQ8/P1u+yNjMg0UrJhkEu6iPTtv
FrzMhhi5v7nMeMHn+SACpdW/Cd2oKCZhWtVk8Nasgeik3RDUpuu6M4RCkum2
tS87eYST7P/RwGO5LbA258P6g/FHU8gGJ15w3dcOuNehfa+wopUT1g3bPZiq
OXdwzi715WBFgmHjGSmxEmJp3RThNvY+zVBzDsrovPqJ6opQKy5DpFvML6ra
JlJxNrrZu1zUHITF3+ymb4H3XXvhLS3qmLG5AMYNOwWabD0liD05lKIJtbBE
0hM6n7l+nZBhnwfLDqlhUfCmDGRM9VzzNsN20UzMlQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jeW/bOQbRTntNzu2jcOhOb48lcDYXBqPfVyQTDch2UrJ1DdISGtNT4I24qQE
GXO240DFJVFISywpfMp5JlbfrqxLvtDTXVB+Jn68nOtr2DwJKc5m/QgiJwPE
+f1pah1jxyvCPEq04rKlRV/UT6UuG0BQbShkkneb8lhNQas17mM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Pg4HFiQXnjv8AwVUsACPwYtiPz4ryiKzL14G4aXEUA0QIXZ4utVCJRn7Tq7Y
5i/PVtaOsZRayyrvyHBIjs04uOPhCaYVJqrLMUUe7BnI6tU/tTocbMSamjME
xYyCWm5kx8CqMgvxYsNBPwAFzBTyPtJ2+hDETdCq7yZ/ZMr7N5dnqtMp4vwt
oENj8+J9GjuBaJZ51ef/nUXVMCBfG+cB8P6wzPu6Z7JESpnUCi3YbQ7SW/mA
w/Ey+h2VhqLMmYJ3wc7ylG/yxRKQDxmpxZKg7tUEbXR2n1yLj4TU4SY7OLpO
TmBgnOr3Z2EA1YP14tJQT54PB3+j8A6gglgkBL5X1mHOl8Cy2cjyPvaPf+el
mtY/uOTLZidOyNSchnzyXm37c2cgs4YKayUHeH/AXk0mA5qnUiYnvybunl1b
8HbfDHGO9Qh9StlSl6773sroQfDKgwbH9/OIqq5mk0ZRBJiTCzcehHIL9XRB
yexXOMkNVm1932pfblOLZcjgX6pc5ADm


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
c8r+iIFMyToA09iq4naZsgnE3NTcH1MRM60uT+r8HvIwrqmeldOYyE+uAQy/
g6XjAZnKom/+l3ksylXhhGT+1J5SBO6kOVo5iRDBVluvsv9v9uUVkr1osaoU
asBjQJN4IsH5KNxy5SJYQZ9ttBgO5ex2dcCdk0PSPgEE99MW1sc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DK8vA8yYsbodAPfgyMbP8WyJ1fNAC4WNOIbLMovAbekq82VnAmBTtlkCAuKx
IgfPNlrWG9rSvHKisPKVWURTWmzjKKi2zb9bOk4EDY95Zur4VEf4Tb8qG1Lp
O51m56TOpfA6SAJgV5sx7wiyMTHoons7PGEHIOmHX9Aq9LY3cWc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4752)
`pragma protect data_block
PGPaxfeh3Ai83IELoRqtF74HnuUGnD3OvlekZRLEuxY4qLxvpkDuUQA9X6KG
xmbNyBBYkafu6ghXcY3e1AoKAPj/et1uo9LsxcyuvjDmm5vUfdf9xqwxFXSW
iI+eDt5e0LKhLt8NBgqZXwtDNdhFhK/Db5LW/T/GIZLk+ivcX1clmDTgUWpS
WEgAo7bImXMww4MR6jJGsG2NUj4kQBuOI5yi1Lf7CbSkxTL1kUcm4BNxaopf
KDyAtNqqsEWXGFLhO+RM1noxYOdrO17KnGrDy91VZZ2I1bX5J3RfucULEBhs
V4L/6a79dESBCMLOLdhxsS85jgOM/rC5tf5lTLnnn27wvD8HZyqRKsTJ5u0N
AFFma4KslLSNq4YZjL15S1V9fZIDRepZo8V06WmzZp/xp2sP0idjRtgOjPbc
3U2CQmL+xobrgsq3jN/BSzLRcZEQZN+CpEfDAZfhjTXj/kTpezTBdEcYSc0m
omP0Kz0YoMmSpCy202Gevx/M3WJKjf4n/lAXHBppap0N/pOt7oBAjZ3zmFUW
3p7If0tSLEBNpvC45NCHK4jhD+/n2okNIDOr/BroSN0Uq8hQpiJ+dYyCth2m
3fC7C7L1+vw/3gg6xpXP3LRb9m0UnnU8N+Kq8JG5yUHxnqeUGuONPtiBQh/5
aoYCXwNGHQHU75tQermffbw3DV6vRGNIk1bhARFIfSfTJuCwoEFX3jcgT44r
VXkEWIm5hhLS8XurYQ8+s9+JTpmhSfIYfHvK4JgBoVtQ+2jQrgRfiWUpPK2B
PrhOZxAZab74whbkYLCAHH1fGDVp1nFofJyOw3S0tr2/vb9hbB9evwy2OOKe
tbTnb0kCVOu4Q7BsxFvlpjCmSxPWa10mlnv8ge43eB0ngfYvMzJ6htaRhh/D
hADlSgX7b566xi4KfeDvG6F1A5svZaw5y7579K9jl8XalMtwK5jcJDuuAn/F
NvEA98BsTCmaPGzWGcbnKt8d5QbdWiM/zTbBuC+Dhx8h9oby50cRgwdzwuiH
1mjg2GP+Ovse5iqlU59I0EQ813u8p/Ey5R3TC775QTMeUHBPgCGcMoyjx7TL
P8XhF4gxzGkDQ+qFT3bWRKm6SdfpKqx4NvD+gwjS+rCjpNIF/rSYk7KVyjAu
ZZhIMi0KM1b/eKkLsosZ4G3gXVKgJ+212YH2vS57BMgjXNWgQqz164xNkN+f
0VSlEDDQVd4SkHHD1GuzwX0cNLhSKQm2KiTAtR4KmjBtLLTooiehAJpQBH3R
ZStaqztxQR/pG+Ls71zggCGXbxJi8wIu/I0n7LXwD2TmaPM1eYUSv+QQwUCQ
AyEmZNDtgTQssIyCtO+thaEO7flK6yK5P7SiZNby5b3uBXJObOIycsweQnef
Z6dmKu87QjhFSRPse7Dmp3RBxcz+1OB4jHLsrFWuan9Z68gLtLgUJrAv6VJO
ebroXzUN8skMo8HuCLjjLFejZdqV9osFIXxc0CnrmtXnUM6Kc8Hsf1EBHOU/
SWydhjfYfRt+qU2DiGDn58Kt/MyY1uDdNKYHDp8pARkCCUZ+iXTn1iCj6CMK
M90kW5agZEykeK+3xItOU530Ud2KxXPyTmpco//2jJQgbll7OnHJ4GjAtfvZ
ljAtxTPnK3NkjNquY9F6lmNmz96ZRRcYTyprfRQUZaAHlT7LTVw8Xa8i+/iV
RV76mxwQf3HSkRaNZwQD8jZENcTkcaSxbpCbszccPJ77VZdRVtGOzgam7RYu
vrbaAANhham6J98IR1x7FWuO03NaKs2Ihgkunbp1nfuJjceBNWC0sn5csiR6
/ewGB48cqI3y40Mtb0aoIxg8DxfeydGbfVVaLC3UjmVttx7wFLSsUIDYYGCm
QGZPwBb263r7mnz5xX3Bu/Pni8PtCXp3daiiltzSw5GX4RnJxgh/0AiwFrcy
SCeLSpWC+U6c2lMZwaatHepU5ih84ER75ET0VjCBw7GGIpnSJF/VqihQgyMv
rdXG+ITggA7UHzkvGP8MwsGDF1LClKESkkxHucQBWRAjpJ6m/Enz+CYUX7YH
RxYWos7USE2WD3QGCqjvWmvfkJCPbxS6Egg43pX+UEZjWzuDh2sd4RMp8/9D
rkn65PygVW6FNHM5VvKkloaXw/zLoNPoWDyu6CNjX782B1Qi6wYZaqfDYRTw
7c0Cd26feX5MauTYzlCDCX6AQaQs+c2GbdNc2Dn1DmaMOkaACxTFElGPSXXs
/N1JJPx0xK+AEs9yN9c3WAT9Fvsc3/ZafO3TU8y2GmOVKPS2YGLL00Y3TOIm
fhfmWipQPIAkTeNZ3MqyhrKBHeSlKlprL6xdDAAk3+HFe8187+ZwlBcgl2Lo
2B+MCkuL2/2tdybTTweq9l6zIIKUm8a6xqtmgv1fZ4YyOPlZjdABDsMz+HL5
0+5SlSSa2MdObuLs2cjYQqcRyf/6PoQMfRdYiP3BpNK/lIqQRCsEN9StkyTf
H1YbgdKCLuinE0fNqxp06VLCPTyPsIE7j6vVuo+ndrbbo9zUvOfOSk1/vVWY
GAy+27O3WzxVnvubxtsf1ubvb5pfjWQpkJbRhmmBZvltWb3JRKIizIw8qEF1
y7yvPY1C0ZedikCG/4phxG46hQAIu7B9v6XStdsx3OKoCQw4QPyw+5IuzJwi
XzHneNuNfqNDEMFL7uhuZAy5bW/CBg6xyTQTkcOS7w/9OVjhwga81MLTjkA+
qJIjXcOIQ9ewy2AsmivqVQ6lAzwD0njImLQqnhL1dfIaol7Y/7dXiKFY7na7
iIRj1RB/twVbuCIbKInA9KyrFzLQy0xR6pvUst5DEBHox60CeOc5JDNEhDFE
g+YWZkXiXEdm6ndpkZ9ZPWZdP7ABwSOBPfEReZ8xtSOn8ysaWyi49AXUe6fX
yyHZLVGNziEGH0XzjxMuU88Ki7NByOv6vO2fWYb7vh7k4Cv2mVK9gIRyV2B4
mwKvTNy9bYKAg3ph6OIRjA7bLGIzbkAjuA3iD3kUmR3/9v23z0jB0u8aNybh
sIt9NUFXWpRBzOn9NvH6mSy9yL2q1nzZT4keMp4Q4WbpyGKSNpBm79RXeHER
uYTjtPO7xmnxO/xLUzD7bYHdB2+TNPKJ5dOeknUtMcAzdqCIzT59jqbwYBsd
v69nxvKknDAwmE04AbHpKOTWbjUSooGTDHe9UZHg2xXgA00HNdGu2LDYqiXd
O/JwwAVxHD3BcJtci54CxDT7wyXinCCd1cNcXMdLFNwZpj19rkerj0d6P+bk
WWfhQmpyePJezEyE+mX1rnewRan4QYvmi9UWRQOOMYU3v/lcRx+vhXx9cqIv
DFHPAghvkEEVMLW7vqm4osD6B/bByeFewlIcDTVZk6C6XbIFHkFgzBvKIgRL
bBodnTecyBYEv/255aTr0BbxFKRsmRYrDQUi5T0uVmWW8jIwKgkzes1KdyMc
5iRetjqp/g55T3j8JTTVGRdT9lUT5IXvrX8tf7Qt+4S4BMv8xOcfdeKWoFyI
jlVOaiLFVXDvgl9OPKUwKC4iOpzOJerxMgTmvLv3XfuS01uqoVrnvsaz78UC
hkEZ+pdxt0CL36M2L89T58aAqxy4tBGbfuDzC6IA5Wen6o1iANjyB0HkTwYG
Cyocw73mRkPvD8bJBthbAK7OZEj86n2kgElQQnS6zPhAcmP46oS1bxGybTxW
dB0txm7taStbFMNzpkwXnyS4lKjed9QDsAI6Q5QEbnIk8dpBPwbtv5AA/0xe
lpGr1impovyHp8gjPEsUI6dXbSiYepsBuL0OUD8xZqY28rAKKsFJYhDkv2Lv
pV3YL72kcC2uqqQDXz5QYftQfN/DKLkkgK4NhdLlMNgUAvaphUpWy6rrXqOr
qAgpABM2aYZp4+rwwdO3pvn5c8rSshN3/Lgjvg59d6HnQfCU7HTWkwUqvXYX
DApEgi0Ocvh8auLXFjcTXSZo4sVIc3PGRjbhoUt5CKTHWrBfDqQ58rFCOCE3
sfDG3mx5uiPDQB5tE2dsxrxl//k10WSJeo7RcjwBXKZgeM53AMQqwiwGM5CH
TH31Fyu+xcTmGQHSq6pCBvnOnhKOVnhFLEgE5/R3ColbZcbEXT8lsx216Ytw
Vs28KQ+fI0Vx6moj9Is4foyhd38R1xeKHH79f4e+/BhpUaDsjycMx/XYzSGe
qyQ86vQ5hJgxcaIBqSKO0QKdoAIDqyN9SxYEs16QUbYiUny/Wu/tugnfXwLH
+NSa7oOu+aVAzzy3SA9jR1a+vibnONlBjkVoYRikL/rTlzUsQdlzbA7bu+F0
gKEzqcUsGEaeoWH4qb+rG0hu4XM6/Q/b2I9NVISmhiPZm4rVeGHKSPAe/m2e
j6A/hEnG6vOt7t7X1srTjiD0qvfj9TVEGAWUO9rOAVEziyfSJV4JyAGDvxtY
+o2tFTrbUMpJJfQKDoWdVm3Lz4j7tobWtpQJQpJGbjfNZxMhpqw3bqNJFTkf
mQiGaLn2cEcM/pfn6UUpg0Vshgj2Dz4Yg+WfqIOBs/3si69ogaH2vXk7M1Rf
hxYBZzuvl7Ea575KGO5i1a0X2Wesr6pVxHi3C9jDkWyBvvuvYFb/FCLz2KD1
rFeTEpEfcGYzVvLQ1WtW1z/x4MW+Bwi+jXmTKLszfthw96r0wIFFKUZi/s4A
lhC3GBV2L3WZi/76AuwikNKGz6dmAh2FI5ntDyNeHEXGXEIFhHGp9UaPWUMw
ZWUBrQntBHlOXJ444x77vABudBxjBhctzxSn8ftwKuQg/slnJG/qKt7cCfBP
N/pDnGNd7S/e54l5zBH3IhhdFJpJTtCpsddOQA/ohK+cwIqmasD1oqhPdASd
Yze7kPRet9eeqljyV5Emyequwi7Nz9QtNBtTiuWObvDWq1mHBm0PNJp8mPda
DSPdsz0sI+HNVEPbgHi/Uat3w0P+GRzB8rmnRjA/gUkhSrs3rSUomBf6auoa
63XjZ/EhvSZfz8NYEPX8HItc28Jx5wyCeml9+B00hzvtuK9PidlRgwV/qBkH
6WEjcrefM8ltYYiLLDhbF634tnmw4R74894zIFg1y0PP8RCU56IBQQ5L/2lC
vkKIR96ZnYNz559VRmzZc3H+8gqhdbRwv8d2bwo3NHqABUIhQKlNbdeZzBaI
qHB5i0kLu/XExkjN//iRho2cwWeeTPLx33XuBth19hp4tXUs8N4BhSBZo3Ov
dexwfcLZiFO+36puVkDO/XpO6QgjGzetWlSc/umoR6Pikz+p2Kmj0VElOKH3
Aen+Lhykga21uKc/i9McRiw3nkeym5BKFCK92No0BlG6F54XNLgGyD8xzjV8
L58FKe9n/aLUogmG4cdftbjjUIeDHtsXRvx++NI6PazIcv+LNbxnyjNwIb7y
w9t8zd1VgohJTJS45vjeZbTjSffnfdZ7shlVKDD5QiA9qtll8xMeTCRg0NYh
h32GFX3L1bNFBZIQK6aijM/Aks3YKJKLsTcV+y7N7MBgzSOvrcNRhZ6WGIc+
qT1JMp+GsJaRcYCb7kfXLkFJlP3QofRkLLIxiBcQ4A9kVUv31F2tPFYIju7p
jQ2h6RqDKSShGFQsQwAt4jNCEVyCYFlLfz7e377by3/NP8ygBpGpfPCMWJHA
qH0MvBrnM4wAwTloxvk9DINn41FC8Iixfs1MBGFncoPrBFp6Nvj4he6vraxI
i7hS5DmiGpf+qpQ0okmEFy2979zuPrisEhhp4GEfK3QrmOT8mbLtmNTN7HN2
yMJskwB7X836Hzz0A5PdyDfugTfv7yVhptP/mcIgCljgijtk3UNWZqJAr5fb
jbpPnK1JTVHy7Qk1Nl9D6gwfweAp4zEhUivj53v0GlGpn/zCvXC56C48cYfW
1ImXJqAL5RvQLYk1K+4o+eoI8PyidsvZKF6+C329Aipzlk5M/eKLda7Miorw
L4M/IXsGP99j1+w2pOvFJQqBZYI8JiZEsb/p8zGR7sdSMAlFVKZast5XgW1c
XMOyFCyQFMxpa+9WMNXuZhWAvKnbRIoM8Qno5YlUdpOGJ3D6tLUQ9aabolk/
ZwVsoIw7PoLxAGiN6Zor+E0gDMaJfbUr8ykA0MRd4La2OeoEV1gGa4OVCB4a
Uc2EzP9rxl6jMfF7vCoxPv+1BvoLljncbrgTYm+VqFRAUOWqcEZiM1Y/TcmK
0KXA0gp5Ly1lKaMMg21z+c7p/ijDBKtm/bzKoJwksqJ9u3/b6v/gRqkm+bDd
i+/orvM18MAcocEHGKqLg5dD+XVvyLfL87vLKC5yx1aLKx/grxNW5m2oOmko
PGjUZcAD4xwKWvkePfUEWL5D/2GXFBeO84V44Q12ezGt6Gf+lStLZaAR2GsU
Fboz3lt1cvnFy2HX82XLeG7nfYhypU3KLbCw

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "cZl3+z0J02TVIcH2La0evC8ZU8jd4Tuna8DsuwukiXDpscNI1u60Qb+Bc10ZOZqqtZ4tU/vmhVv+F9Ysjn63+ggxQTfKs2i+Kg923+dlDx5ogYUMnCsiUjNQFT2K681kKnmkEcWzfeDuIZUQfL3te9+bwCurNMuLZIKNyzpeL6wfIikv5UkJ883l6EkRUqZ6PRXqY8A29Rf0Y0sxDVqm7tAncOf6le4GAj9AGwyD1to/d2GA3C0n3HUjWeRyLDaht/e+WfruCZ3LEZ/pc+OOm4CE0vn28r1+E1CHKaGaRT99Rtq4llzP0GTpEeJOM7TJIxsQEbLRzggN5GOzpRDEu6+x1kJKWn2ulP0Va8+xfuIqB2o7qOj9jvGX1Xy+1IOnQVc0r3HO9la43q31yJJzsQWgd+oU57DNdEhHl00ymj4NwM+w4B0jSBOFuxltbxqldbjtl4YGk8m159fsr9tQpxA/704MBgxt0SDl/tPqVGjbmMixEzFVUSxfqIfT8/RjU7xjhMRApyH+EZ3pwAmAxQxwWYLPmFaoXcRifFcDKAJBbISpZAMt3+hbKx6zhGzqVwi3LmZ05ihs6e09orwHVjWj834BtxVJoLiI+G+Kd7UnWmezNEQIO1ITvS8TdRer975ylDt49FHep1LwOXU50x6YDk1492y/ADxeDPkQXk/pNjv6FfxZB+CmE/h/H8/DHoi9mRyux7MLsOEXCDQrT3JiOk2+SRXSN23oweiA2RMI7JIayJ6smQ4SisXYLkX6jrN5n8FfuuJBUDDmK9CsDCAzGKcMMjPSC4Oe4TBYn7/7IZN0ZWeJmOglfyqBIAYdM55qr2rvT96RwsbqnSGxUC5/4Yi3RBedF5K52KNG5rw1393399kdbEKYKHz4MwugnRIyeW9K+w8Wom2hEpuo1e6SfpFS7IAuC98iJnPb2SxHNEPPFHpEf0bTxea9H4qQJ2MBRtQlcYEnfBc/LeyRyQRL1QNlX3Pde/2e51MwMT9SlUgqS+y4q41BK7PxRIwo"
`endif