// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CSI7kjkm/sGAlZ6GF0RFXFzFzDCaiYafLfSK1Qpl9Ft0nf75kR09JyaN0vSw
2t/3hkuWcDW9jJ7hJUjzF/6rRwgul+t8Rftpvgd15vV2601o6XWyqFpat4e1
2tlvSz/niqFaP+gT7aGLptxskjgaXgtAHyy0RiGxRYB+s43LpC/YZeq8QsHC
Co8ENyWPFR1hhhnQ+BotFYiHxJUptngZkztRGmUqilMEdyGdeLOfyX+3Sker
P8Xm4e8paeEoanWZcvUwHAjHfTqjRFyhiyZ0ZvCvrW0/UZIBA3+EmTJfBA5o
kQlYN4Kj6a36PkenQcOt2dKme34zM+hdQaMRMlhLeg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dKqwxiRYH+s36szidjac7rgix4ikobvYOlTJfKHU5cxFSFZsC0gV8B18OtSM
wfDUeElrB/t/Kx3aP+Sp2adWx8Q1mf4ioSqrl6L8MXMzA1GfVIVx2puNOteQ
Whrq5rTTp/Lt11L9V+I+6mMD8x9tr7sUmAMfbZZBzWkaWwsdcSrvVWOQxJtX
QF91DVws50HDNGn8mJdCqYIeHB4Yoha8u/fdjqBywMiywqwBYAcKq1PavwmZ
zdYfKEv97cNkbM+hRR/10DoAzkt+RDlYMZqrfTd2hoaVQ39BlgP2ig/iFdSN
DQlsrHY0wfDSNC8tbUKP69M2n9DskaS+wcvfT1ohsA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Bq/eXF4xJbCLQAyAYWAZBlgnJ1HtertaNlBLtr1CVT/XjZPS+DveJt9JNN/Y
BsTyiVPfN3BsUU9GHrS6SEHov8cYhknWLmKdAmKvFJYuwd1aps57zR+88Ge2
R2gCnBn0OkpaKoWcxr/ApGZS+QaQ/On0PCg8VAg32svkV7AIFL1D9iE77YWV
ze8dI5Zo6lPmR/Ry2pMGi4WPUdrld6AH5eLOL2AVMPpeoYSLt99mYCjt+ury
q8SpRO8wXMVvB/d94WSqlwXPcG4pUSL3Ek8tksdV90Y1LUHBNla5j+sZQ3Ap
MQkfkzaLjogpORciEgZwHVkhBdeemRm6I06f/QQUhw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UqMsB4fIobygZaEoTSnEP9eKK4sWG86bLmxL4tu45JWefaBCpqPss2l5+dHu
raMd/LBm8wt4hX8RDf6QhEIPs1WWR2KM8OX9glqIev9AkJgdFNbNUBpFCYc9
+mAZDh6TSGJ+jgHEErdOtaEZxdaIcI+w5npeOdemLnMzZUTH6d0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
lcZo+uNou+7ldlgigZV1rIz2hWZkapVeR1qo9gPOqPB2i9FzA92wKn0OYvn+
F1mgdiS5Igmx6HOYwbhixkrxW8F/k/6pYB2YDZ0mYdXk+SLL9EWHBEezusXk
6dc/wRwwzNX/M6frHkocf8v7AUlZ2lLzhs1gLakBZzbIjNyRQPIs50tdaJ1V
vn/cIRBn/k6/LB2D3584mV31VrbaKeiFYaov4o0I1s3SZ5eAeQUZ5VKjMjSQ
IudsuckA6BhITywnvw1iaGN3nJOYcux0bvlTvOt/1reB72BHC8Bgj48jSqvf
ma043IthvER76ck2XY//4amyLCub+MEvCN7aggTlm6rQpoRcy6Zf5WkEgyof
iVJeAw/ZifGpDbu6ksQu7VQJhxoCSMjyYufgvqJm6wINoNRln9VeevdnfVDV
w3pr6PJTvXczBsYgpbC4FcqErUZ4JdsuQniuS2VUmgZt2w4FFOs69xbWTv8I
KB8YWOjqIeAQuC9fuD0brW8V+nlH++UX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qyr276ZvhagLdmix+XCkro0vdX89KA3+7+y317edhZWY10r602cGvCvSrIeg
40Rv8nYAjmKTLfPuqvWZEZ9Q6KF8qs0eBUzrtgS8zEEcWuqYVunvy9BSMoUV
C1vAoW8Tc5QOlctGeYEdqVdqeqggBWoMwFLL8Y5sT1bxraR+R/U=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nqrkJLF8n3fBR7B95Kfn3BQdzE2v0U4Ee8VMOJF3/AK+KWtJTCDVRF9mK2Fr
DGP+6WE2DhWH4fOCHuVY9eut3OrHOMyDvzvQa0ytueBOXrH+Yst7yQDge3MK
aDKphHxyDEmtz1c7td4Db7G6/8kwYIPc8uFRrWuc/Bt9360OBFE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8848)
`pragma protect data_block
trVVGGTVzAKa0IZFgDZyAT62gbkKNa8Pjz8uG4JhOrQIPdV7i2BVfXLh5FWO
QgrzFZgxUmxnTOseHBRzKLSQZ6zdmMWIygu7fuWfC4gK/Kx1aC+Xll5c1hCs
CnUGoeuWmSqfuq0ZRT2Zji1BzbynbtINM8kbT41x3HEl6dtSYzMYbx0CEUu/
iAI2kgXO3vEau3A9OWugI5JnoBPqz8PlWbAW/U6NVL2oGz3BwlN2A2zAo8ci
ik56tUfRXcqVMzl9+RDzzTxaobEIWjTmRRRSq2orfDouar9Lm+2H9cOo/Mpm
UGmaZ9dH7EedKPBYSiaT8Oqw2ji42zpx6de0tGJtJ6soip10/S2eDTUrwvVe
48OkJ8zyn/TlD2vrpkoeSuBMwbr4oxuTRD3pIqfULsm5MIGRBdeCyttXDEAI
kjFPFOfwR/QjZjPMOXRMbHJ7kExV2XKmvIrdz+/jyXfhjIjst6dRXAFwQZY3
+x07BdtOHikABUtCSzDOJB9SYwCQzEHG5NTPGQwZx3LEMwvaZ5y07WWU7XJA
l94jTEh7+wwB9Yampvp+U86BLjHZKwFuDhmtRnIr/XG6xizUjpsfdnUC95pt
j19dWcJHTzWIT1bMcgtuak0UYp63NhRDWLIPrq8gO/7ixeOYHTJH0MpBHi+N
C203gulfDBFtLZD7uY4rBFhkEM/hgzaa7IKL2SBr1+LJwi9astCxvoK7uKkp
fcGl2SjSXzb1Rn0xwxRfdqRHmDq12WDEkreq0uLBhJ0ur9XqIVcC6ESo7a/F
isTxFykqUWrrq2tvB8gho/Rok2iBq0/mRoVsSkU+wMbWXIbsAaxwSb3L9kDz
TELx3mQgL7W1v2iJeFiDAJCi2tS2AzHp4J/ZqTyMFBLftUg4u9wiNiuGzP5e
LfFDbWxvDsGI96Q8p05eOpiM+Sd4lJJK/hAH0Chutssf9Dv9Bl/P5s8/DJvL
DorW5qjC7h64MQhq2dLDJUMSmTj8PbwfdJqfK5A9TIS25pH/5yhOQL87Wq74
x+EvQ6q7D49uUUN/yTu4HXMn+XuuMUHJwixV/ghX5XYVKTPERkwtkbt9Nk00
e8/8PDjxnwnwyW/axHI1uvytjklNFjUsQouF0Au9yPhdrsrApgN1qIj1cWta
uW8Rd6TWwwsA+NNNTy40vjQ5M6E6hNgkDTreP14WZDFwHCLGoUWfmNv4+fXh
w+hm6hWRte3msgWKGCtOI1hRsmkwJFbPreTQmWRiXW+QuCRx2RrfBCaoiaXQ
E8ZUJr2I4rfgq2VrPV/mqndejGT3h0V178AY4+LhKUFAh7jeVtNaGTfdapKW
WbMulErfWqNmHQwWX6I9AKKprhNUWXmmeYUTDLEX6vEiAzOZVGT2lGP8Z4Jc
EhgbtPCbo2jz8h752Ucc4aplkaDc/aBqFNjK8jJmqRGdSlCAryoqTCoOfxwj
GttrgWnJZ8vRt/u9MV5DMVPtxWrtuvxRTIQLQ4wsYycK6oNuCaKpEpmJwpcp
69Jmfjv5iuEf7m2Mfa+MVti67ki5jXQAoEYYUcv0CTfLDOj+oKg0OaXSJJoZ
Ovt17DE37IDplSU5O/mwFEEabnGYx7WOpHzDxovysfeB7ZivU83cEYwk8j/2
FIjfjnw2NCgwKyT3PwhWOGs4wxLCKOkkId5x4/SoQcnL3yHvKBeVFiw6LbgH
ZiGHKhOybrYJlZqOKxeAmYtHiL2L+voEOgkGJU/VtNSDgPYBSUeiq7h17HCV
IwTNSKPLDyLtckA6la5Z9cAxVII3ghZaJUcUajNnEQ6V7dX5JGUU8g/p9bhk
WicYBXUaQO1ip93B8EqDMlNomt9aK9l1rfeE44ZlT4i4IKyMPUjZP8qDeoWg
vCWzI++MbhldojPGDMsNlYEJ5lvtPU+X0bGo46mO9Adya6O5svdO0AJMnp3r
x1DZfUZfDjKGtGUu0doYBJCryVCFjulA7BNiEFJ1U27LjbhzHR2x64TXN7YN
vlJQEGt4XjM2EFAHSGTrdjmqRSVw5WfQokzqhtf3UpopYjYw6C87/g4/3E92
tMxjEtmQbhmPp8nsRDAsnyRIrMrhj+Nl/1I/8BXPp6eW/FB0WI92tjjb0eB7
7z6kbmBAjxzMNXFw6EGG81DG9MvBuRlPVMIYgF5bb6LRY30XF5dkiIyjcgtr
tjoAsvZsBEekNcsQ7uSDBj2HVT5QL31mHyrI9ek8/2kYbYwIXw1KoNZpNIDY
kTqn1EM+e6hDL0GU9BIQexr3XfsRvZON1FnwIniPkujyyrFmRU839VwF4v5D
H7TEkFK4a4hTl+aj/HWnO3ygZLUr4y3/Kgjsd4BOSQsHLFhta/MRyrOUSG+D
UW3Vir0Lw448A8VpuVYG3SUxS0/FRcR3l1UMMaawNHnTSg9Hrnyk7iyUU+m+
uefkVlEs/mbXp+v6sJbXohCIeBj3fnSMIH2DNWOczdiAyKuQNgSCYzllbsXg
9qw7vHUnrTAkwvzwPBfUiXgcITQ6Lva/+hHtwSFxKOsvQ62ByvBeU89sBa8P
0Rz4AdjZB2LxKPbvTeNW5KC8Fyt7WdwX2A87RnpsQkCL+bcTpE7Tqkcx8ZSg
8+eDMsxNgpFguf4NJLigmmb6e3e8fZv6P/wHNzPrWU/f9yNpR0RouhAl/xqB
IA3+rsZNSCO662nyO1zu4GeRXIcEb6Wr4CrbR5ITYxWPT6PY8nSi2V8opvOM
hVtgCyeWoAEReI5XZTRHKf/UVJbREFoEPe8SlYxQvCYKJ01x9yf+LflBy+Wn
do6EI//yC8JDqMQJsaDQOWlWgXEhJs4pAB0qqy0dsFNqNFQyHyVYHGCns9NY
dYR6uLH1jTT/oMa9zJqg/Fw6WmIxrweYrI2QMixjKF5ECvf3z03ecTfW5ZNi
cJV5ASl2xGE6OOhOik9f4TeESuselZAD59FJR+/+Wkn95M9epXJpGQF/YKAS
K1JHgvQ+4sE9W1RUoxvzQF54zi8ENZDQB9Tmsbk3r5iDA/M0+Qxxlst4s8Sf
n9Nt6dUVonqizKUjOqdxpxt7frn8hVT7yQSa2gI2FQhY/pO6805tDoqwJt4C
jGRT4AJJoPn3BmJEWl7PkD0R51Uj0Ybxn8LYUFLEILZIAhzY6KTNnCG85q72
67hzbkx3gGAUUXbtdMeYwvxeWf7y+A5WgE5wf6UEGDXq122CzbNchtUGjlZD
fMxMBZBREe8+4tHTX5J96+SWEQ7R/ff1Amy+wmxp7KP6gbsd9kZKB/pp54IN
mOEEA9zGq1ON0ABsdJpGytZCeHt/oCNEqRgJGtMZHSAPmGiPVLQcyRErZlfH
5KGmEQTLVBLh6IMtrc8SmLNqKZgX7RRYrKRbmXxIT79nqAKtc8LbmfQNsSTn
lFOONVfH8WvLUsllgiMSsBNe1moGorc8KLRX714lYvdmcmg/yFxqZ6In/3Q2
EUWM2G5b1zZqGEfD8z44FqdlS+ftPpa+eQT9Eo2vpILRDAJTEflC649EkwPZ
Gl3Jthj9H7z24oPeSlEf8aTfTmcv22agd+pj+LlEWgmsTgD0ISq0pH8zUmbX
YF+ZLXoMUuah16GLidAAphpArSLKX7sHTW+7JVlGqvf++MY0F/0DG/yzJ7wu
lUEf3jgX0JV10ZdWLk9F+0TmP7XKFpJVI8TtOwqPV/b2U8SsGhIV15rD4UbB
7WVoxwhDL0Yl2wkov+mlPihSl/x+P5QQW/mkLVSkZKzpfUnyPPCSF/5lN84h
mWo5TuDH19hMwemsgWIoeUWI5YyJ98nKsC80VANM596q3iNr+DXRep3XENXC
u94RZenPJy+C8AKByG4ncdE8t8+NPEbMf/9xcdLLaZqcsJMhM00L7OXtkrTL
9XsSHwnEKBlNsHOsmW5tKluxGygyXpA1HyIEuES8c7hcLSH/rfg2lJF3yHUY
idnR3GOP+uvMo1HfsUx6W/HMCcBukK6mSh++ECECmEGdgCqnKAqEpnMQq3uv
2JjnlSavvcYnAI4xkUrRuPtw1+nlTz/1nnsN8Ug1uduClER7XzBisoUa+qZY
+gcyBe1WAv4zmTm/+wIj4WJ/pIlgB1rfalV2TSZcSdHSFllBrHhQDEp2WJKK
yib94UALgyNyUXYNuymFzJVoqgc9vRDDsPSCH7FZKA89ohWnd/qdKZFr5DZ1
cEtCelKrcFp65b96b+wOsDgtSIhbeDAPYIcQOURgdeXA/UDagc5ju7cB2ssd
tKbdfqixCUbu7qfXpKuLPnSJragBZ1wAZFY6z//eibDZp1trius1qpz5Z29H
6wgPp1YuqHw36i/OrRmdYe1HnpMO+SI4LntjSLgIwK1AzSS3MjOn3ZMFedfq
TA9ifywFcFfCXviXg/USusSfnW8LNJkZ0LuZjzh7Jg1RCtj3xsC4EkK2oU5H
Jcqu+eqlqvVwavx3b5Gx9tuaPdgtuWdwBmLrZPxvwB7FgWHjV9aF+ETPHR+P
28ZwzFnLAh5JJJly5/7U+QTVjwik6M+nUrvDwp00sH1XYRsMhFiTFx8Ii08q
zt5OvJvU/u4KYuZz7ndPF+uDHWjtD0ZizC5iGm3JP8sJIAZV9Hpnn7K04ah4
jC5q4PBXr+Xfxy3982Sh3jxbPZg4BHbnC77BdfPF25WexVxagEuRymJedH7F
wvPmJpqoWZmIv/R+4E06DevmpbbJot8cUtRPBCjdKcV7V9nK7VLIa/V+2BQi
mQes1hJQy2UFft+4iziLWGN3Qw23IDHrj+RZ71U56xWC5QrEr4JDeAkQFDUH
27/WwDE7jbVGVSOXUQchesC3mZNihdySLRNHJC3Rx0KmApTbSlYj6dMVeTnk
Wf2L95IpBow0i0QRLACxhgaD1IeC0FxCg1PrMv4lnC4RLWsHtq9r4f6Dg6MW
DgAIHcx+95G1LZ7ip3AYohdI7IjjiMw7VAh5RQzeFSq9EC2Ody46s5PRUgzK
VxXycLf/D5m6cRPCthJw5O0LHy5en/8C13XYyRH+pUNGKRZYsTFucxxCxmm3
YdRWPnXq/EJ/+J+y0a3ICyrQr4cFmek1GMpAppO3BT1uyYdP9vKJRj6WDUBM
ys/jK+hVUFVWq+bFEitYrnAtrs1o5y+OR72Su3OzpsgXmZmtA62n5G+l0aQz
lxx/hznvVBsXOPfCwTnQZIVqW440/3OulI8/rmD2b1odveN7YgloMnDPjZos
O28GyQ7KX3X78EAq2D59Yx/HmxEsxye7jewcmgcNGS3mnI0Phxlc+SlS4X1L
yT89pLqqQ0+6NNpH6r/165Mo0UsJlsmesZT1gBJnBzsg4jlYEFsnVKATHZfp
OehnVm40/hYopFsUIqB1H8GPkWsg36L6Qz9UmgZfVNlyD+TQ6bGfNyJs1EGj
XVQpJb9ERit2bhCD1uDhmgiRivsuz9/r1YjPdNAtUe/BnO5WminxCfSXM1gl
+CwinPUhWYbEhoyfz2Zzb7OfMZ0GfwcYrphimG+oMYgVXtY1aFt3QAM7wFg2
sMrDjPf4d4SIkZVjpMibegHhTmvL8+ntKv0TJFQwK5l+5sPAI5IU2vhKlNgR
n6rYXULOggFY+NUZJxPvELfxpP7FAOdsQefjUNBrCAWFrcqVTFg08M3B3erL
SH/N7yiNTxiqAuyNppmiXEM5W5bWyQ0iH89MeaokEWVN34gnHe7folrK3bjc
94vaItzDHiXn7CgqSfiRRifoN0k1cRAGTRgg2hhDXq34pY+A5wV5YMASvw7R
uyZkFmpQCDvEPFVs1yWcvytzhSV3Jwl7A5zJ3iMppzhmAmPT5Mtx9/Q1Cnoz
hX8q0J/A4gen3IAjYQM8mruJGjZgtGbSNnKC+9SbscVTF79xMMLJ1c3RBusN
wXKuniEmnE/mwaeUJKEiKImWFWRGTCGsnGtkno4YdpG/wGrenKSFeCiIDJEc
Cj5SskC9Ni3dt95LagXKh+uLJKMVzFvukJBbs+jzZozrICFaTY0lq1aAqNb3
BIFrMcZ569yrL4FHGbIZyrOGbK9Ufe+y/EWC52wLRvvAVz+jzS2oUZhNfYLo
jQ62BRyR+EZUQb0ZLkrNdJOuXcrCmYRZuWiGR6wT6fi8dEUPfz3kHQA+v5aT
F4qi1AR2ZjvTfoTVSH/rlYVwmEai7ggI4PN4pHNP7kAAomddo6wYmbxWzSbP
zEVLrSJSqQ3IfOTGOTtsm1HpTv0Sou7/WFahZlhOXKeit3Zj5EwXsqqBNoOG
FFjMQhPvuOQhb3DBrkKpwXFrNO56XMLBZV7nTmLBedyzoC4Bl8mkh4/wdSBa
4ba1wbT8Vss2wNYp8DjPJZJLRUZPWRVxDG3HFDnK01bl+gB0Hj3MmsBrMeBc
maPmlb+r8kMlOTyhBDLyLhh76mF8PY2xpR3s/XZaccFKFzPcsXK3o1BjPyao
w5mW/vcV1j9Kiyjvt8I87Ry5Yp5d4a8qe8vwxo5WGEnjYBh71hnwDb4uu5B2
IcZ/p/2u3/K2ci1LWdFQ5Zxz2TpuZ7cehjysQCGzaKXQ73OX6tSq/XqLii1w
DlOjMJBHLa9HbKhfcaGyWdfVxKIJc5Nxwz5/2AcKJQsl3NLKj5VtFqM5cF/D
jBODBC+2ychNTmaU3ZJwTbJwccapBJCmSaaAT52gqVw2jvWA4IEBlvLv2TXb
Oh6V97gFF3oUIZjU6r6NqTppDMRbXi7iqiNHGbiboi8R8aAAxY8LkSMHyX/r
V0kmWdMHjtSro5vt9RkrFwoHbKGEetVjoyIE5MgmsJSpQVdr0x2CD2+e6Sc9
UR/+QH0D9KEX+qjIcb5lW65FQocmiPzn3WXtXn8wc5QAsu6aLbzLJUXVU21/
VBCdlx5LZnHsp6EFdgDoO6MF5dqVsro24iUXES7/6uWj0l9OMLLbnrj0mu5q
Q5j31E2UtzXSFGOAgXZRkdjdqqme50E2EFTBagHCBCn+vsMxCugBkZoO3fWe
fsNPS1GZCnAJ4cbgrecExRMQzGZMvo/CmPp0vAf40QZpWWXlI/biq3jyAnYN
jRebR/jUDrqJ7R+gTsEIKC73IrZ++8eeG2FTFjZjXvL/rM/XJk8dLGZWEH34
mHTadd06O27vttt6G/mZp6RP3JtWFVJgLmD6bdo+988Xfj4HRikF7jpbwV6/
zvXKdCNzuoDbno5Nat3wDCzanytk240KHiKGLzJ2JvKxbi7Qrdy3vSG/zWZC
u3gQyNZ7A+agWgvtgL5fGIczTIC9JSr+cnqPfWUohVf2wFDnuNaURjr7HJ+t
v74dF3VqoDak7BJ7PtEDjsK4yDAh7Vtx8YVwTrkszy2HeiQeeTSAQ1VJ3mi8
m0GHlYJiP/GXu9ZhEZyc2ZmCmJS6Qed1RZj0YEVbfgiwiwQE9D6sxr+B1mo6
dLdNFZRlJZN3imH2eLQ1wJF2wKXT4RQrVWFeS2vp/QUKNIHIBnA1qtGSxB+D
Yc1qogBNVLJN1qRZRDmr1mOze4rLaDFLyOUEgFVhBG1Q/HW6ROct9ubmMFuW
DKXG1wDQfPBJKRAG/QhXfkA/2ns5QPp0nQ69PDwwzIufZv0Jnr4A5nG+mjeX
BAh5rKjyVKkWc4qUjevKl6aN0z3vgHdEUUuT3PwOQIOpmKZoddPDcGAP2Umg
Hz929hFvVdchl7qZl6oSUiUh3FNqAVNedL+klaep1EMSGb9W8ZUCRIG+mNhP
IpAXPHdBUD69YuQgQKyhq1hKAX94ywgK5sofx0EuzFA/Q8ixeEv+sidG6472
FMq0SOd62m8RS0QLMN0S0ZbDD41S5te8AHJ8nrc4riXb7j7os/aNZBPtEJiY
zBSjTyNH4vgAoX6zwI2PfmwpBL7Q7HiPrdbObL63Ptgr2pnvME2TlX5FQsXi
kmTscWIMH7OQofLzE3Ta/jYvq6pHf/hW5GBIpMwRZ+rb56lMo2n4KD1EXqAJ
kGRfyv6FVR+EXDMVBCc60ctD1McZReU/M4LLbTd2bb/EnOfJ7qPNCIFq2UMC
kaBRhThr4a6CLxQoG30aMw/4vAyxc9AYu/pxPN1rGpcZNO1uZqCbnnTShdAE
Q4yzrhSSIJvXMuunrH0veG8vl60dT1BuBb/TF9jMuNDv2din9OhJDeXhcCjz
gDccnQmJsDUpCJh4L0uVkmvgsJI9f/e2bVoyVESSQhuMyb4Npc70YpI1ENQh
EkoFYMqxIn8KxAMKjjD8tpd5OXGHSAq5HDzIBgCZafNMbwyTKa/eCPdYvqaY
e2v6ArhQZOwuSrcG52ZbOKcOtfhPdqJc5AZFDEM3Cyce77Auq6IRAr6Ficnw
CEUpcR0EC5wbPQ7BbpDr43OZhe+AU9NZpWRL9P90jWQLQCsm/46Ap30ZHWGT
KIW2rbGhFzqVKb7lZv3w4ZecdghvN4OPS529be/lFrSPFG6xye9HWvDDFSi/
i/txlw/lYg22sBkgpiiV8WIZu0uU6Z43+Yp9QpJonr0cCfOInkAaYxjvd6RB
I5P2D2JDU6lEjunYCY2JtWlbsDgwN4MKHYPZQ2YG43iuDHGusqWJwnXQ1134
S+pQBAN/kSB5S6gcokHBCuU3/qzbfxbSzGyWAg2qg6/5qkkLUNVDE1UkwBza
xE0o6h7LhNfJ/+vMHDUCCM1ZAHTzX8Yn39XldIaXeaF7AuQGllmG21FCc8WE
5t9zJY6WxvpPIB39PNPJR86qb2PI0pX+Gk3ZKxqAd3fff2H/3WNvJLIt9Stt
UHXIB0alfsu7XAtsfihBGPyvYvNWYl+LhQvU3YIB+cP/93DV40F0Xy8iXJjl
E7kLOdhIP0sfU9ZGeayjx6ir7oeI7z4C/iG3W6UlspEcypn/KuGVyq5Cjfgb
F2LnRsCOqc/fhsmjgCkORDFnREvIjJp2M7pjHqx70bQROKWyn65U/DqREceZ
uakUKxVDGrp9hGXIdKosDZ1s/J8F/mgpTdMu4wlxkdnNXgVr/8QXgXHLVYI1
Jhvgki+Tia6D/MPmOTaWYHLuvG699JVl4M2oOV5AkhL7LR0OwKlp/EkJfbxr
nZRtZedxbbSISvB2/2yj7AdXheRqHIU5VpyaWMHEH9Gn+4/ruDdElC1HD4Lc
rVBy4s1Tu/HRestz1nGaKMlJ2CiaP4jsRzn+agCtiNPSJ8C/h13E4JSKS2Ov
DY87mrgOXHL31GOMXMANFweHWPUA0YvC9kCExtL/2ICVMQ/dOb33q+FWN5z4
R9slHdQe7KBhBYEZZzOoLnYhuXpEMnG61qnHyUX6KLaX+1jEArp4e54QBgJC
qivZmjEWSWNa/X5GJsaud8+8l77hWlC+s/IErMyWaFK11ONL4PGr+5eLZx8S
tR7tBhuBbbtYM4lUshixu/en9KMmSp9LWWBiWXEt9T+sOw3ItYQ4yOoG0ik9
z8YNzRd/t5TF4n34HRf6JzAWHwooq8KWic22MF7pHdbjIjimdfLtskKZ/zYB
Z6W6CMsiAoUFULv3+KUBGngAMqWsEHiE/BLtEe4XecIJWzWYMsM9/v1N/BDU
1IWEK5ckAbX+kAh4qvAKBGS5kbJM10FPALpnxGlrYlh9rnCWk7qKUikYbZzx
+EcfMVlzHHJWM859NLadft1Ll1ZHkeYjIK/QRO/+xP5fW9Dk/NR/OzBSYlvy
J2STtVYA3zNjiPobn71tezmb+AfzJCT93PfTey6q9njPCQ6lQxNYzRtTpWXN
RDOlqtwed315rDzcv9Il3WBObxVsj9tBTURoaj9aJ+KrHiuMS/flBuKDrOyb
1P2c/SYTFde1r6OIE5hGwK4Voa/BRzFZdpc52xizEf1XZM26sUb4tMI19uFT
Glpz4UmW4Jy+rHTv3WQAKi7vURDuhCQ1+dbOkbW5fdJFMOFd2hvI2iFBdQm6
JGd7F2NqU3i9ttTlNAgODbtBQgKCtmgQVz/JAulX29EhoQQ/ECySOkI3+gFl
EcucO6DRYX4NfpxIqQMmM1BOalzCrDGuC4z2ewMRq1tiSt3SEMBG53SaeepQ
0TL4tQpKwO0SEw2I/e2Hnd+1IUqeOZ9YhAOmULXPciZaOrhSSkXyGdotDtHZ
ORCGgHkrDm8R/+hQM0M6tnookrwmZY+hb+Wdk6b6mqGvDVQLalAi1EfA5axY
B02Vu3EsPOwwjZMsAve4dXLvaBSsZ3b3lwnu2AHbaYRo0VNxNEOtRB4XHgnu
LjpUn+Wx+fP7ehH2Q/gO37dnGGMkbX7j5ZK9s6MzsRh54gNetiJWefNYUb9H
NQawLGhVcG3rDevei7t9Z65rFobChiUAEmmTvTJ/+tMdtpnmMWDTgECxbKA5
VsIoW+TexzOKICbhqv54l6CET6VJrSzHGzdn4jm9aT+Q0zsTzvHbsI4rX/Ya
02YEQSXxuM5bWHXCoA0C7WXoYXvJh6SdqIuRreUTANQRVY2hwcIirtCuI+Um
pCwbJlQeE9sYmUxshgOTuu3zFYFqNjwQ5zsqcEg63JdvOYAJGfO0Hhv8cwHI
4U4Y+27K3oZeOMadXvdxNN8nOa7pNiTmHEtWF8644i3XD483pyn1pXisu7FU
NeiH2XUfxAgXW2U6ooidcdQnE65RYrwGMaofhiijcBAGM4+WgUYPKcaMzexJ
H6Edp/ajzrbYP1d5LUPzvv2smZIga6GlvzTyg1RmN2zn27SxSX1b5GXqwvN5
K9hTHi92j1K1ZiV729DfjWIT+8TAxniciBiSmzPVKoVJ8M16TH9d9syu6K4K
HwLnuubb+hLVHxCMIUOG/AiPbIpIER0OwB7cGCxg31BmDpMmjiGicDQO8csy
SEBf/xutInsr2z9UJ6P6rzgfWCPN61ppI3Rs54SflcSD0AaN2OW65loP4+oD
mtR8ulQZUrqDobwlyoBFhYkvBGWhe6e2B+aiFtMSuw1vkCju3Y1ZGQ2BVvQD
v02b54ij3z4zLlHOobxOmJBknGoidsYJioRqWCoI7BI8RKsqba73FcuUW415
NdOzY9Ewrxe6sFNYpuTxt0CK/rhEAKU0blJHN+88Wdz7yb/E4oLtQKbAlg/f
T+JhmWsjhFTUvmOsugsDYo/oT4aHr08thk+tPdOZ035RR3u9AnBIqvRCPs1K
yyor4ClvIxNeJiXWypG3VLq4+vhfU7t9i3BOWykEKVuo+EU14LpwawIlVRPb
ZUYfi04Kik5MVRGKb7UYEMIY8BMm/QhvDqK8s1newXSoPhgM3ywbjHTTbscj
RJP5oc+2Xj4u1cFy0XBWfVpzXCC+U3CPLu6yMoJCfq6xhKpl/CnTRHG4zIBe
/c59OlJVtk6jUniAqj0goDUgMxchBNFwhw28BzEjasyZIaSpmp/jqHccIFpj
imnhxwuUhm7HqN2LqbGrQ/Sqj5tzDVNbvbGWCPWvCK6WnY8YeFrXsBIbdwRA
Xjah8LJc5qEZwTM+sWIEAO7ZqewEaa8ToN7bCtDb8lpk+x/QIPhAcN0/lIM/
K3GXxPywXB26FyCcsHQJTeY6yZgKC6U+afFL5xbnBFAz+nmaqOUtVWjPid1l
1CUW+OBt0Og8vLoOyvTZW9fSu3Fac4dO78Gd269YYEwYNdN8kqkn/axdJDVP
KaMUaWXsh2Z61sPyNYtGYVcdl86+r41NmnU41BSXRdvN+IAiIydpXvJ8CvaF
H7czV6Btq8lnkPFF8S7RGXhTALedHXmAIESJqLhuWTNaOy0mrGI09lUDAXQ6
+YdvgiSDewF5gilUiQAQEE5w6zhtjSznF86m1RKzv2BYgS01dXtCkaZQ9cNo
EWHkJDra69c2uXvwawwUh0mct5ofCGgPE7SnO4qX/bUuTgtoW7DmmfNMkI+d
jJg6+e1ZxA4fXk+RUJ3GLDI4iuhsrnkq+vyVGhdKsUpCmIwoLgsmnPf9rAI7
4/qUrT/CTpFiFqYnHvDEoYfOrmxVA/lbiQWSFw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "cZl3+z0J02TVIcH2La0evC8ZU8jd4Tuna8DsuwukiXDpscNI1u60Qb+Bc10ZOZqqtZ4tU/vmhVv+F9Ysjn63+ggxQTfKs2i+Kg923+dlDx5ogYUMnCsiUjNQFT2K681kKnmkEcWzfeDuIZUQfL3te9+bwCurNMuLZIKNyzpeL6wfIikv5UkJ883l6EkRUqZ6PRXqY8A29Rf0Y0sxDVqm7tAncOf6le4GAj9AGwyD1tpNBeE/em/SLvKqNhmy1u6waEA8IC/hNZvuzgjSRKe8WyZFfUr2pX0eW4ucAnRAcD3g4lQAxgmArhSTLz124ikSUlyZyKPG4Isqg8QW+qZTgeRnVrMnqIqNAgjWByHLPgjY8cAMf3ltcPgO3+sL3CET4cNwxx8JZM1SMdnf9p4L0Fk9ZlPFS+gsmTROLW1lcfquRSgQAcaPK4m3oqXgFFTqwrfgUac1D5Bmkw2gIRtoAfmlDmUpECoP4cVA0f/ScnwUIBLFSqVRDmZLj2qaTg+jBapGdwDyWFTKw2vmM5+mHXrJreEeWQZYDL6UR7aUF/wlIX6E8gPf5Np/xlDk1Fvl9mLe5teBv19bDiNS8oD6eQEaIbOnMGSt0LEmXYZxTpNEDgrBK5hHqR7peine0+5Ib/UifgHsw1Y96FZXPUr1Z5Th9ZId0OVQgpPYRb0fLoO2D9fIKI1RsLvAimDsAqlDtgLcloGChuLXhHQrsax0RjgBpBVXJ3fNykuvdtHXptA/qtmqnUtpz/JpvKvhdABLeUxEOioV0jhe1F15nDykJ/kierIC+rMV4NdS/JXwJZ+4pnHUT7uYaE8hof8U3te+pF/e2cPlvlGZlKX5KnJ1b9gfmXalPn0+f9JD7xlmGkp13QNmgPm/jJAromwT8qxMmPwpiawO/XPYDEY+2Q33vTXnkEocPHDKpGQt0Pm23vN9WYx3nOdjUD3nxbTQhEEzPyNAMhEq/kslWwLZckLU0VATyeIGKFbXoQrI3IoynI0+xvXFZGkRXL7BiBxH8ONG"
`endif