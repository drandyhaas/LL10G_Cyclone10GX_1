// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
r7CR0zuh533of29GUzkam7DJMAWUiY6vEYJTkla0goOgifV6JZmeDk0xUNL4
BL8LfkP9hlaBY3AuVTnbhAoy2vJylbP4xVpF+u0HtU4HB+t+QVnd0Ds2NGxu
ELqBE5ka72rDm9cP/VfNCKGkbr6VvLhPFgg62xzD9ivNjvWMfHh9GpalanZu
YETZSGbPWk9D+m94rqhj9URTdU4DGpntrP1g3gS3YmJIol8YhDOL1Km09C/u
vv7BE+C96zcrFFh9vcC2qCrxF7kal7culuUU4eRtkeNSNuBoLG+F9pW/Vesw
4kVvb5n5tyzYBmrxYkMxQ+ovP5pAlnraIn/tZulVgQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L2S+Ic4n5uvTu9o1hPjABbmnhluIzKGkKn7E1lhNrwj117fcfNCU+RKT0DnG
qB8oe3LzD2DXgnP0U1sbmUN+hAGm5HcW6fngvHocXNcxNlc65Cz8RzCd9iIx
bAlMX+Nr8nAZWjkyhVxSfmBkcaHgjv9GI7YIjzfz7oKmD3ZrLfrzf0JV562D
8MwmdbfXGI/EfdPkztIann6CI0q0hHfCOWeO5l6WCqWgpN58ps04ymmT625a
i7hTnWLi1j2m4JClCE0QjKI61Cd7RO40LnGrJVAAVzYYALksTs46zx1E3CE9
Y/K/eqEv5yjxDoMRDAELK8ViBzyr1tB3oQq3v5EnWA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bV4LV3dDtuOg8IvjD/bmFJqDT3Zbl+M3k1v0uylEQmBVJgVR4vkl5sAOxspq
HC4Agd/NZdkPbAhEJmfNPS4Se190wn9BcT3JRKQAHrcngXx+bK6KlkbZjsEO
S3QFFR+aWk1/t2FR6WvMER//XgKg/kRd+ZFoR18iGQqF7TJ5qHjETzlqqWoS
uNOIdcNcfmjY3o3nzzhIR6D8S936JQrqVC9W8p4wEr4IPu8U6zc3oidNEE6Q
hjnnZAJt9aLITOHtSJ28YMtRKO1vwrFfWeXh55REq1rEmjtKFsfBp1ipFhhN
p3E7b10JXW6KiNtoNK32+BKc9UgrF1eiqcueHF0ksw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jrCMBjMek3YLoGAIeTdM2TyxMPMFrinPpFlK0zwQnoLWtw4UgXgI/97QGT39
aCFTNT03HQlLmooctAIFJYb90HIRQAOdhknZBmYEGj3kLuARczx3G2Ax2Xku
q8OjtUj+cvLp2tBz8rr2X/euOsvH9rVD3up34Hbo/hRkQ2b2pqw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ZopKYpjdRt+31yCWARkyt1sHLuC8/OXPQpzAllh1x35h8AUIWMlWt4K+E6r+
s02v7OkBylEKaUlwuHpbzAMcjf2rKzssWryUduljlmoNqBhTlIkqulj37ER0
PBJ2k+MCCaIZzfOFecY7IR/rXzaBHyiITTpO0hYNia03mNU/ypEPD6RLYf59
5Mvra4CHi/9lWN3ZMMJgEUb4Wh8o2QfIJ7opbwiqJLZr5ttb6UbubCrA8Yw4
nRLX3gBwNJvchLIF4Heuq2LpMUOGUusUDiSYILha1eByDIjFLoW3QnTp6v6h
H4so0CdPZiFQhu61Jq4ROwXEo5Vx0rjmPmgOuWYvX/VW40U2F2hhoYiCoeNu
g578wOo1sqoqeHUumGOuYoylCWaESu7+ZL2hIEZVNEcHdbB/XKlHZNOAB6f1
t7lRampdIkZdPDmUDVZIjBr9ss3vYGGGzVMfVbQN0eLswwiQ6XoiV3uqKQMY
Frv88XQQv2gipenDmMMTpPuvEKIoVS5i


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KI5H013EfYO0Gq4Mw/FTF6+tclxLN8w5XAOwlWGpi4oyY2r32zx2j3ls2rGL
cFebnxkE/UsDGIAEnEYTH+jvm2kKVUPLN+LVCo79QCln2LVsVht7Taz9+nIL
X2RjFlcgZIwLcLskRjIYncxvdTICURZY4+Pbc+DYF5Kgt7XQE1o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p5rQFJmJ1IxlhaVr6vJKVm2NaTCsuu9koLT0MSKfwYV4bHusRZiCT3l8xcBh
6KgB07xz+ET44pSM6F1xdImJGSDnT86VnfRODTF6UwOnQPCFvPU9etT1UKuh
uSSI87JMx8mTCs0Ks35aRxovEIdDeBHydtfAlVS+9r0DpPgt2cc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 58096)
`pragma protect data_block
cQ7/leiOopgT6fkLrryt/p9j41ScHALIVK45ANNojhRpkkyOwvGxdyl+RNt9
uy9rHsFEFrWApZ3DZwbTzGrWK+PGDqz6pDO4sxB8X0oZLjEQAQmgAq+o0jw9
BKa682QvOHOYk12J5ivmjYnXH7jlPjI7wKJunzzwN8CnClxQl0D0KBS5/UX5
pef5yGCVTIAXPMdxp6P46hKsAy+io0KEoJSpfjTBwqidugWD3E/9ixyERtq0
RmtmR4HqOIc5FYbL+aZ1oXehuIpXR1pghXmuDCNuE4VUxF5VkfKw+dmkofb/
SDrZw31AACYkVJz9nCsFSBRTnUpENhiHEGWeZGqhYAfRDH6DWmi7jNXAns1o
vLWzz5PsDyWOBsBqcXhkbTGzi+ktMhi4t1dyUAUoB3Io3opPYZ/wlU/uP8f9
rBVytfdzJQ5I4gh8NtJYovU9fYsMTz2ggqeg4p8fXo7rkHsQGylJ4nd/VGuJ
guFAJGq4RJw2UznOzBVOfm9iJSXAvoSdonBNepkeWGhudYKE34yErCT7H7aP
3zJ1Iel6J4EM6+zIzBq9e0obCVwcBO0Sx2/hf4xyP0TAbQ67PKQG7tawdCG4
QHRUdu6jm0JWAUx/w2xVtEV84pU+d3QLSg8M3y/R+KhTkT9sr+lbgV2u5QS1
DEj32IT1wZxM9N/pF2gxguUMpVJhjUQPaAWNAasIaBpdNJFBN79LvRpVxkHg
MWawnO8mXprF386NV/h9v2MX99jWsWpzmtn+/Fj+VGqJT5n2Ezo26Q9a/a7F
VYvKeZdOuA8Vb4nBmlxHIbNkY/RyeLiynOKUK+2EN4ZlKlS2i8ElYh4C2KUB
x0YFeWJUKu4jHCikYrBVCf8uy53QYFfa3kWySWsslG4d03TacnfFYSMAPDQs
2OUrHPMk/fQk/viX/BY4zA6rvCYHxk1uUzsX9XJ+QA3Xtc/fHE2VaoFreYjU
RcY1q+k6Wt3zvza84CLrlzM2O3fYpUwDPpZDRbDTuy6zOts7/9o8vEoaQVoJ
cF7t4wQ6CXBKjRTSQHvQiv2GHELCpSnyVX+paNafyy3uitIjg5tW0zy3CV8P
ciK8eh3Dsu+c4Sfa0SqoQbN5/ZDTFwe2xK0zKUgcd9aJRL9E73oLjVJMvb1h
GwgscQlpp5DjJXZ3YJSM4ad4jyUYiYXPKOk+MeZFpwA7JamdhI0nvibS2kXw
j6sdU9wSC/7jr+wDqHTp9/kJKZvVUsT1YzY6kc5N4cOO/r62H/BJrfqo3bVw
U5eGFksgH0OHJQp+DlePwqEHFaq8EDjddHc4Niq/JlpKTR7nhMiic0vV8i/B
9AjANtoRIIIrACoyDFv81y7/7uKTbBPs5bQruPUaBZPaYc+bNqi+OCE6pzxu
1v7mho0z9PCP8rL9dal1rCEUyf6oMTMrwN+RH7PFE67y7qje9iyyFxs6+dyW
v8CoaN/4EHER9P8U1BIygbnCFCVKq7vbWnNyWWI2J5F4utIQeAYa9VvAFiwR
9UzPwibgxUEiFHD/rvcFlgcIc2likfSBF7Dt2/fzsDwbZbvjdduhf5BYOZtC
qtOOKfJlFB4s0+XqyCP7Ae6mG3qfTRrPqasrPfJIMvspuBaF4GhBtFkgOT6v
1UUbZg48c/PUlWwuaAje8chqiZarYSAVM4yWUKWcLs7Wq+KxMchpbtwSY4+i
pOUIbOU3DGfImaVBDe4d4zrNQZfmfU8hkk2FGlggSDBkM82wVP7vLS7NcsSd
A67RQDqEQCUHhEOfD2TDkSg454HvCdLq+ZvFT84ANRYXVjaAI18kKrZPyjne
T8AozGUpj6/1iC9HBqcYiYN/XTCRB2lgDd+wdil3QN+kGeAr3ITdjE3YnWle
RoHRIACwPaIykIeso+bf+0PCKQ3g9SdghBa3TbImRWcua+UUY7nrfhjdSe79
OKApjo1EWGseKWkGhty4vnChnfesR9AQkWp7EDdgrJDdcP4OqIwu3VOAtxSL
9LgpCsK1Lj/N+IfLPTQiXvUIumGphLJnsG078oWUeDsTedEgB60JKzgjpTGE
FQ8juHh9OtZxcIHJGcmFwgVxLxyH4vRpk4xKfS+X10zuYQ/FUUGJCq/fOZqx
5P3YKhFQN4vdgpFMr543Yvy1QbAhKkRdhL4Wq/sUOQcH5BsFTkgnYS3CEYra
0Fz7/ztWnT/HPBzbLkx5Ec6JhxcM8D1+lhQ7SN/PjfMKEexyG+2d3nhlUTTS
jC4gHUDaBo2BLLOOEehQrA1289G6XwHXFfmDV1PcNwPuvCIKth3NAQncOfYS
5snGDbnGaB8Is/w5vzTcKgv7RnhqhGUxvmyvXwliRRSdNOSOiu/kpWMuwDzC
wIrnXUHtZcrBca2AqC9m05apuK2yM/E5UPAahoIn3hJVEk9Ktg6NPPcCj1ke
sGnhg5WPs1NLC40Io3jXgUGeT3N+iLxysuWKofHIUqM6yqW8rgmzdDPm8HlW
szRsldcTmDdppjJ0ePiFYfAsDxIZcwcsgVb9MmCH21+buOM7GBEQu1FSQH/j
PJGwSGSfH4IVszVpYUCzJVnmicsJQhU9K2K9QtMYeWqXCDsZwkegY4Amk8o+
OCAGKBv+Rf934h/Er1rxn7B56+Vm+gyxJA8egxPFY4gz6GxVRJE6+wSTJZ8x
2WYMGSsEDiOBVpCJqnI2Nzl8AVQdaFj0osuUQWiLndGigh+efdhtl7FK0R0b
tlG+wxJ8GZK71woo6heoT/N2aQLYAC1EnhoJ6IhoEy0daLZoEmZG4/D3d7fa
yqAb5c7STeZohQxw6Cg5a1jPUCSOwWMKER6ViUR5TpN73442sLrGXx2vTf4U
ilMcHKfd7eVfMDjyH9GagDq8xqe5nolczWvHQnKcqXWtHE5YfosZs9vIKXC3
eFB63unmz3zMbCXLAfXT7xTBQJJbgpagN/c/gFR50eT/TdTvA+BIkB8eFZWf
WLXaOmZnt8AzuYuBhktle8jFPSjL9MVqvXjJ3AKMsi811FDDXTUSA40GmRbV
xQU0mwGGq1CVJ3q9jZ0sqbusosEXNTZAFHTGRbRkMbDoafHUl0gdLhyMKlxs
SnnoDT0tiWFMFm4WBpfl+Pcx9xJz5KFCxIcPoDFO2OYbviHQN2WNUKQL4CPn
DyZnv/rqjp0oDfie+mOM9fGkOalJlmRyvWAsWJZUcU9pISp+DQqYzvkTLMju
RpktedqbuBnMEwXKACDHN5iyBsI/tZIHMt+vMsaKsAUNkA4nilmWMccEisSN
TN1weGcIE1ma8/EsjAP4bjgWZiRRBrRrw542f5DCZMujqzcB7PfQaNcq1N8i
+U/mRUk9RGh2XMWzwnUwGXdTveVE9tcUVgI54pcxSPxNd23wt1Vz9IMiEupW
NqI+qbMLBcjHfrP9D1jYwgFEOh5bYaR31XvzvgcerLyWorQqnYHCJsfIriIp
XgNtAB7kYajasnkgy0EMQmSPnG3owI2pnMUFxkELpKiJTAhlYe5KGRDTFAu9
wua2qCyTB1KMWL1EnwX8tW203OUq2I/LGb6GFsvfGkZh5BZLbMr+PbJpgWbQ
wEDXS9OkT3AlyM4GBvnmjGO31rv5ceKGf2h2hR0vworYU1DcwP7Ok3iY/yh2
XaW80H3DIotx4D4QtvjoSACxqMZLfu8Cmj6CbJLSpkCfNB8otUtCfWhejNNf
Zs/lvcq8YZ6T2Zm07PFFcSo4HuHiq/uVBVAqbCCVK9AGTmwofCzUSYL2rWia
8x3qfOdbtDm3wY/FonZH3CbNzcovuFN6rFa9DIKOdPOP9dEn/3NXnZ9HFPgy
Xph8ptZ1T8xTvT8hsnd88Fcp4NV2Laz6baHT8h+IbmI0tkaHDQa/3EVkXWFQ
xBGyOQikM6fQLvDOgacYLSSfgxMILgWdRIXK2yQTMqRms7YSrHcm6MvHUjGH
X1XmOOacTK3jGqmnbkV1DyuxlI64wCw7fKHo+vnz2VRgMzbd9Rt5enSLw33O
mKpqNE36/XC2WThyMwCMMXT0ltVub27Dd/i4o30vnqwp/E3s87/X91X8OZ+L
0O3ZJeTBsdaL0lqEqsimQSZrdWKICB9skQ9cDPyDjIa/jXeypZHvh+DRCJVu
Aw3YQOIaLERT4/HztuuB/SXzUJgfYjeTXPM048o64c9ltaHEU7ghygIM/+/+
Fepql1qzMq7lJhJQ8/G0MLzTfz2OSmnG3IVmQWoQRAUY3isGvYk67zBiC6Td
K5sxn4OiR13fKFO6LZPrHHt1Mmx7vxifxKhR/fSqDUkvvFcabnbf7ISAjd/l
TEaBrNeG8zSQ/OQ9rxWu/qyNA9GYd7woXAtYAzPh4l8oQBhPgj1P09JHmusv
eX5KNwN4+hdAQHs5klw3QWrrkI1K8S+lk2tYPBbsQY7P3f7WKrj3aJqkcrHm
u4j+VTB8UqMO+uECSbiH/jGaSt8kUJOP82LUZmXFvVDTAXs8s2xylMay75Bo
r2nYv68V/0teASCaaj99N9fp5ZBGgS2mK7wiVkbwG9XKggUvU3umV9tJdVl+
T7aB74lH4cE8waWqJgaYF78txXVgApI6CLNuGC+w0Upc5U/El8ML7RZUImp4
MiI6E75IAWBbXMowbtoKlo/kJrMc/7qyilrMZ2eMzDMnTQwVUjQbvgS+0GDG
rD7B39jpCdZiwJcQHa0s9kZ2QVOxiT84yP3GUyKdBSC1W+YuGWAPdBPAV52P
AInX6fHZAqXetRgf7rMmxx/w/Qap27OuDXp4q6S/CIStSa2vcqrQcnqv9y9B
0sbFazGWVIDc2rkpPC4MIZy3nBYVgqIJHMpFTeJBadWNQ+HElYE7s4xKeGmZ
00Uuy7432hxktreUTBDmyvS4Spv7zG50v//u/CIVYN+w+fXfo40abjlnUK3b
M22prSymgM59mSl+JpYpoiJa0G432Qe9jPIgXXINymvIRGo34OI3/qYqqe6p
5KU9HWq8ewTrcrXih9koSE02sJpdR0AIYZ+LVNaK7HEY0eFt7Hysi4sbKDhi
vut7bYBxWKmxQ3cvkDOoW9aECDZbend1WcYCdsPTFHstxIJ5DXoHlEddCG0B
S3xE+HGTMM5F6McyKHWQCFwCvJlFuionNgtVUG+wY1PJ69Br7Znls1Yd0MPP
xishbs1hl3wnDnZ9wpwV5zRkBdmKI46vG/rToLmFZMCzcLJp3TMSAJ4+lIiu
+8NWMMTBtFxnlVqBP4NkvUdpz7kj95z5/g3OVQqWFBmJ5Tiz9EXcE6n0Ia6s
kFkQM5EJIyWNhbNSLyGFn8Ov6N4jsjLMPIXoxoN8JFydIjDGwtpDBE4xpMuR
l797JrsWnXX+pCEtvQ16nDSeh3f2ft+Eqc049AceJ7nSt/inSpOAGa0LARaC
ZpFzSa48ZJ9zjxyv9TpXAfRkV/8gjoWVdDj1C9Q9Tw0Ckp54If2OcN+2NJh5
vjBPm2MR25C9SsuQFaYwftvtgRZ24iaHpCqxZbliCAwaR1ifBNBxPz8O/4hA
nSvGvr/1Fxixey/RFWUS5SE2EZiflFHfn/id0KAdB23yOT9wYgFSsGV3JA+U
dGAnVS3g0/wj+WhFPW5CjeRyR8rCdcUDF/bHDtCJC6f/WWG0t+gqo6+zGDWW
3BBqlrI+AHy6UvhJjXMI2IJnqpRECcO1q6rsLazloQDEZbqK9PTQllGtUeJb
LmDmEr3B/u72GBS+RoaBvYJl3EWlX2bgo1VACLIQI4NTJjhUKYJePY/vU/S9
qAUWv7m8sSSVbtAGn/hsUjA0KHS3cVkXyapzfqMmD1jUCzDf1NeVAh71GQgd
YanpZcn5xRyjbyz4bRsjbJ0X77jRqu+91CiGSUiwwanRu7t4Zeny3ENZwU+8
LYag/LAzpS8cUpx8fodh3ZUKsJDvr4ZhxWR4yY8udrFZvlMf5tN80ucbHbRY
QYoZCCu2wzO49psgJRzHPZ2eX0khzJKV22JYizeATCl7ql0OykhLXnApbZbQ
nL0GiA78fvAfP6/66T3bv6UpbSCaXrzc4zjAfaPKbc/UlscY6/dYkPtSIf1b
GKmHbJmWUL3c1x6qsEJ4Y7GKX7EAHqxcI9nVb1q+UImzroUs6tsxUI6RhGDo
TP+yJBtm4P6LQrhULUPT8xobSJH7JtoXdM81sMADoCbzBXZ4wgPhYzu7gEox
9zJ7o+lEeN5qEMnaaw9ZMM7rH7G2U7xASJTKLtSoq42Ic0NtpDqm7wj7AK3O
Mn0gKTqgWlVkcN72Og0u+1m31X2Rvto1ZJxijxX4d3kZUk+RvvU9WSq+b9Th
H3ikljZIIUpkOTwY8jGr8QQGJgPML1+AohJTzo8CgnKmyLWqY0s7of9Rb40b
umHrgLZuGS5hxgJTIyEKyQKnBrPaQD2cQ1OI/h+krfksP4oC4qnqDn8mgcSb
Sx5eHbB01awWzMpjBBYw3ULTilmjexnlnGXidePo2xwIwgCGfqV2yoAC2ZHB
TjbQyeKTe0i3EOZSTFO0s/6byGIP6AdcpZ3bkcVGa/i0zLYBUGfdCJAQPkNb
o74sKKWBl3r9lAgpeXxMHMIwrrsOhXMw72QOiwGhZTg4KcUwuqMJozgFtiLv
deBwpXz2CmWEwosK4vPaSN9HSGfBiDSc6Mfe3a/ZzamKBJ9QQXPXwa+B3ojd
ewXTMU+6Ju5md4mYnDeeiK5VT3z85mywHS01R1u6jaIUGRJJlcMZITm97tzM
W+5DN4WEI1es6ZE9NY0M90kKvybQmbycCRSq95NtmhsGFBwipTVijgxpOJD2
9EG/cv1gZ2OI10WzROT6GfiX+hG2+sp/RnnkFyZ0vApm2xE2e6BeYqYIlO8n
91tjXmn4r2uytQ0rxKZS68olx+Hf6SCUdPyuNqoxM/NGwrxarQ139yrmLgFD
Qb9VuFzZMO21lKgQx6TNed8+Cseybz+VAsc7B5e7OOojjjrg+l8aBl7bFUsX
PqT7TRQKWHNLEOyH7VlFYhf/RmV585vnSXoUoFoAGwN6nKr4dk3NmfcJ5jSM
eqV29UdyGS7TML/LJ9z609SokU2ALgHFgNRTSENfXP5tHYybmrnQMjcJrYCh
/1Cm7fNjod7CZezpOmhg+iHnX8FqsgfZ/9/lJ+xx0LkmMWeF4fJU1o7IPxOd
LEdoKDjPDD6ptGy0faYQoyTgRWzUrzOUptNyv25pywl73t4gheXGOTIKOT16
rZUcS3Ulx9YYR/ZEvpZaSmIfWB4mFmERgzsPUnjCh/5vRlfdHmfSBV7acQ1O
zgrZmf6GvMF9v7qW2TP9SIQ5kDqNzxeNybyd2w3r+HAzltZxfi3DFpZrQZeo
EzQxDFixrRfdS6TDiDksRE//jUKEum9Whg1pOaLmeSgEuCsfxMPtqW3Chc8a
kPPZSJHyGJE3MCaxmnOOFe754y6RfRMmrrOUQESUyQqGjxhuq2GgcMvuFOUo
3bM+n+yPPObbFYNb4LH9Hm3LSTv8O67/O27hvfV3KbjTCDZcXEum9LVHCWaF
QCc2pGo9u5a4Rsq0BNFlwuDyZY4x2rZ6uoRd5YeAJywMbpeF97QBBLT1krsx
iwN4DaJxxexTjRV/AHEr/+aHPbTYPNN5syzxioDdkn/3MmfKjJlaVPX/z9a1
JogNjrZVK/yRbvy5MiaOm7lsrjT350D8nS8wbIE/XC617tdTqKkHDQPA6tKa
MqEUFFWe+kyOHhTFRw7yoylfNJCrUFSzMvd7r2YrNaDFEVtY5LxkXunYk4q+
w9EDDhiLZehVzdTPNhmhcJWxsMW4oYA0CbS56SoYWON1aDp/IATZh510VG8w
JnGSc0moVbhBcOWCpDnwFKlGct5f7UZPrSrDrKBQK4YHb6HxkGuNww+1//+C
BiKxLuojM8NvmrlMKGRG4QMGHm7RuKyi2SDKlpQSlKJ10QIZk35ol8TIkICi
1WH/z0PFwiYQoo0nRTo2InTAR0flCjX1Bdxu+571fUMbtK72A1Vg2Msa2T9t
pTgvbDE/bzFtFNoIT2fpgOWnpp+eD/0ALclRga8u9cfA+5jr91zMEL1zWQk3
p82NxV+X8djp4lY/t9D9LefR4MGlD0JRwNY0W8UeD2ZP7XTEgZsXxg89xdHy
dHP9RmrYxpwK087Sx9z6qpGh2L1ONiwT8YtqJFVa77IbFLT7YyYVu7T9lOMx
g40hWw4BVxjKBr0WbDIGxFSvvHV4mPkveYKs7sgV9mrZzEC7/p8AOf0mI0rf
uDFN+xOf6/qJ+nn0AF28XbQQ9Wfz+VAbb7Y7iRHF+g1f25xVt+YRpRkrjuHq
J9iVBv2q9eF8koYGCjYsKFTmW06Lb4Ajp3YyM+lnp0Qe/QmskVwJu3oysXPF
8Dtq4XnA/MLkC3blI85EXRsXODZHyMeER9bS3d5BZshsIrFwepLkZK2r499a
cQRooMCb+XdyHCzTYvSCI5ptC5zkI32YcOYTalwSEXihhvYWxnGBYcwbtT1+
I4Rq77R7yUH9ytfK2TwQD6caZ0B1QKZWZ4MZgBtm73a2lMLcW46pO/1VArLT
o+zRR3MsBPHm2VGtsexOrUUue6rlK6Od7ef1+xTTB1ffe8e52YrivKRhfvmR
3IFE8AZZABTUs5ZraOvDwXrMhlFZoWn9ERy3UMQmHpY2eMl3yQrGz3LBsZS6
8YaMVlPp4W+J+oIRtzj9GpOBpSb1A/IoJDPUwMIjSq+9H1WElaPbAXNImBBf
7y/BGT7KlbMt9bxrWZsem+tvRqEzkgX07xTXLZGlb9CjDPlJxnjux083wW0d
ixNrxtNtEetBsmi6YxItSNxMthoObWGiX+uXqL5rFyLaY4Xpef3J+WJUFSEe
U6uDKOBG7t38dbxNvdxHBcamIBAYV28+sVgPKLtKPlVx98XmkO4O9SjzDq/C
QqFhUfZDY8p9gXSNMgIRiCAVqt3C0Q6Kvmcv7DVZ/T6WVeWffKrxrr5DWtAe
+zZbjLCVsjL7sdEDNBk95v8IT7ltyNWfslOFfiNxA2q3Wjr83wiQ1BaL/ZNs
b17mle4FHaPm8ZfRzkiHsT+jRnu5yGUXZFKMbbDBXZ5aO9KkKVYrXlZxCf/h
ltKPFSFpQVrFEjA6sqNr/bvcHAV8xLfs6Eqlln/K57GgJtgQJPAuOyULFu7e
Je+NlbL98yfcC5/58CKJoGg/jclvfVIZb3VEG6EHncJTkyROKq6P6f6YXUkq
wjCz2QkCXeSS2HHK+idgJOND8pF1EoACG2BvBnoC+hwzqR+vgqO1R0nlwy/A
Icm7dld/ey/zyDbKEPWmWRCRGSgVQiDql355DB+3ZYcQySLU6/Rx5Tg0BhVK
a9AEcAToFne/8T8WBYBVKVBYcVzVd7qiiztkLdUwATGOHxfZwKAM06Ml3VIp
+jsszzxKXM8vemiEDstfqkz4qpoY+O8JEFuAuhloHgBBWNawGiygb7d093Ue
Nyw5dMlsnUUeO5SJvQOVrSYHk4UNF338xmVAeIKuPJEA93gE3Gnax0wDieun
Q6trm8WObXW1yo7e5uFQiFYk9anDHiqRbQ7knY3KBJcoOL4VZPbZa04fjdFm
uQswYnL/2QQu70w3q2UwkFBc5EYST2Ka57VKX/N8hfY1hJEM0ashkpCBTeGt
gxS6LSNVaqE1BvJpf9LoEdiG3mHutQzyHggTvWHWbOvuaEFTvJdZv+Lo3Cuz
BwmnJMC2nuHS5RaTV6pSxyshY0J+H/SeygJvKHYE02B08LftAJbT9wCPI6gF
aqAele56ChgT/RCh5GDz6Cu96yHvB/mxFYbVV4Ld8Gb/o3SSkvH4Zp8c93+M
TsvqsUOX8rXmHKrAG9/OP0ALXD6dkePGl21GZtDhArP7CYRsSVAtO90hoXFF
R5DLdw7f5hh8D4HvctYB0h68iQFsNeJY15wkSh0FUV8JUoF/n0QuUzVJ7UNS
hMCh+5/zmVuKszpsipA9ehtjUrBvsSc19/llUA0PGA1N3oStREEA014AJQdF
7+8yZBdn6txQZQhsT3+nSyGbEqwa0gIKDUx8yQIXnphfQhOSmj7jbYv9cx9l
DA7WC/4fytnVyFiRbHxLXs/uBKXOGFHBsb28VeCBc/h3UahPJpy1X8B1OuDl
IlhKGx2Cn/qE4hPlYqDB7EH6YkWWTx8yQ+KRACRBL20fZHw+VdcNV88lslR2
nnbn2tp9S6lqZ5YGDYMumm5YufnZKMCvtEs9T9BX2M/K8DV7aFfXsFYFjhcf
qNTFwu+920Qv4nx85Fz+ShlGhG+8bBbhA9rCNJOvtLH+olastBbNx/Lfqqwk
0S2jYavbWDxqEEnPgKM6dxDbzpjTz929cJh+Af2Ln7Ko/EWzgIA8ek790zQS
Q/R02J9bEb4SgMAPquO9TfNFvciLQVzFVw2UUg0uRWcHOJG/0inyMLzUEeFX
0AFjRyAX9VD/nnEErV5GSkg3bfTj/GfSUsKIv+wN3UeWS+aH/yAc365f+eBg
aodrFA9ciYJPH3Tvkw1ChOiFc5Qi1wnFB5fPFaJhM3ZzzwMY/NxCd4N0soP8
HcU+2K487RcxcaxXCX1zNBetSo+qFvhnUYFXSNUaaVazbLl/FOGqe/xRuKei
v35v4dpVWWk4ArBiFZc5Y8WmlpDslTj09flGhgubEl4H3644CkuQ33VNRv54
z11PXqOgli+sg3cARwFl02nO1BlqoazUp/u9H3Ptrb3tCyJ3BHqL6ny48pGI
HANk3hsGtidQOO09TjpkamAw0vsr+kpcZjyqNLR96ya12xJuc4zoEKqNgQdi
IXvjLjt4+0axz9JO86NBD5HhzzBH6aZUexmlN63tuw3wlePkX8//inXQJqFw
IQhKHO2iYxZCD517TgRLh40nILyovrIw4wftKpjcqIFMbn19HitTDdwGHDZe
TxJjDNKFsTiHoCSumZ+3qnH6XnKuaq1w9h/Z4qSN+8sNMhYaSI2WeUTu0r0y
xiz93wXX5dCIDknHMDFth+mmQAEZzHha/Fabt7IVRN0gokuvtXeEAi4SXmwo
PD6IBAwceHMja6D+nrR42dNaDFuLuG9LAFuQrrR/f2+ysw2q/P2Ky52Wn6n8
f99SsiwQFQarPpmqNjPW5WzrpETxAGTQQP5GyK09mahwK0kkLP5F7/mznGZy
KBZcr75Dm7De60l9wiA/dTUl8nOKxc/fnuOkrH0OoU7bJEqjNUp+tCcc4DLf
aUZBPua2yipIRn7go4ksrCvArvkjirCw/5yLjNjoLHSgON+I10F7iaEQg5Pr
WsCe24tw8Z8VVgdkDlY2zDH2RzBo7NlcOA1XCHxsoBWEEj7fM0kHcW4ZsUb2
LUuOA7zx/FISFAdniEZLcwwcN00KAkBf/6FQ74aXKQVFd419vKyxWb5i2dgV
HVzDfX9zgt0cSfa9ciVCDJxXBumU8ET9zmkz1QslbUxdfLjRUxG5hC+vttK6
hz684Yv87l18aCRrrsSEGdsgZUp3XhKF2hd29DBEHxfAOJ11Rp5JuVbVF2J/
wyX3HO2aZmvSzIKGL4RozuhzeMddX2WSqd2PFJB0GD4g/h+2sHVN0MfA7tyF
GYx18p2GLAx7hPiwHT5SytxX0qpOzFSnNYIc17k3BScFdvRYVeAzvFBKc5Mb
HDj94BXSxxd/oBtiszfAB1wpsb6LR3KNruEGPURebsqsWvKDZD5uOcg7SiOB
ticWgGBXt/olIKpwgxWAh+zmIdH5zTPd1JK+o0ih+h1ebKuJ2p9ZGZdZO5Sk
rjVvkwmj+O+TBAcxEeCGQlOpeunRpx7N3P/7FeT4vT/IyowftUqf0R4R+v/W
7KEjA5SWlW8cQv7kNKynfcHnaUHZwsGlV1+vs8HF6GAcmTT4PP55nqEp+DQA
1l1UAFO8xW+miJ60BnAzpRRmb4WYwsr51+mWWP0fHTr4VoY7SlpelkUnmthL
1aZwAXk5sEqVsq09k7DcF4nlTFsqwJ/QGccbwml9tzkarV3U0VhYU+6Lw1im
Vy+AOJcH/5gAdAeKFXRwhLGoKBCzffUKZlsI7Bq+20hmGWnsM7BLgMlO4MEW
7vCOstz4RQlL/uOufM2Eva5vnzQfLY18A2/n8MTBbuLPvI+5zi+ldKtk3oXv
Y/wi924wie1y547LABXYBWMp5MxBKDzWV3OHO5jkS1cFliu5MMQKCw4972m2
b0TowOhie3L5ulBHrlyMskBvCrgqv+WqGJray08qOCkBMzfjBf4uzURMLCBm
XzVhNDuhzXx82WtE4MR7bxRM9Lz95k8EsQI2pGdenKtKZ8a/EP3M/oMEu0kT
S1XMiYF1S9mWwjs9AEMTv123I18yVWGaNICUruS1vSKj3iQBk5Y301ZGTIAU
xQL2PP1O+OMsYnfoou73ESs0lRcmbwfnZsuNT5yvj45qdOj0FHMjRKBnn4ns
Mc7qCca4BAEn89voQOgkkfWFI50v65oEdVN8jX1Om4hb2Y/SzS2dCFhM/r0i
6wUtlPBpgU/azmmmj3JymfDedRvMxx2o/haAFN2ldMSS8o7dHXEKYf40inhS
XHTYlpFWDDZl+TIdpC7z+GCY3ZPbMqJdHzsuCzR50UIHd7kr3qMZEqMIfpyM
9tBg1e+5MwW+xQDp0OyPhJIgSyjxLsKgcMDVyWW3iI7mPWUE8unvnMNQrulQ
cxODX+vk3s7IZODGkQ6rzmBoeAh6afIniYeuR2FpdV/+Zislro3Oq1Jr5i4L
Nc4vJ3aloRwqJm1xXRxh7ilzTu/Q0HsmGA7I4jDqeg8M7TfaoVjTkuvdoxmj
ZThl7kTgNiZmO/8F/MA1/K1F+ToXQI2gWDY0NQMgN9c69XGEJzauIeU26ApS
5UiRIj9qHia6aLegpqi7SphSD/TvpwHic5CxiBa/x92R0QtW6shplaEmszki
h1PnXFUe8OuyOusj9cRPZALwo7YoIhEbJq0FcNCjZ3fpVjnKPvFgPJfzlbd3
SGUj5E1u+BjWzcJ6vZ/nejNCs1FVV5yfriEaMzcWJYLlR4o/z90Ikwt6Cebk
2Mi6iHp1Ce5R9maQ66gLif/vinXcx+z/ZC/pSqxM4m5NpT8lf8rhfqjm0FOI
Wj2pJ2VEbWadRogwOMT4632nlsbSSFfqvS6pJ1hBDmiIewR4bZ/+v4vQAtRE
8dT+h6HaCRfIRFiNESbRz+CQ3euU0O8KikBxuZiWYulQSufm7+4R/0ux0UVN
T7HG2/2G5PnRoU8RaHELvq16g2BOTovyVsuuOP7pVcX4a7s52fTAyra30rLR
97joNd8EK96tahqQw6uu9JyVfeqb43wQNKC3/fDBHGfX5RQ+S0EZ/2KkYhqI
NdY5AH8xR51jviRXpDO9/ugK6GFBuR4dj/HLjjExrx2n3MRhEevl4nYczFDl
nLsh6Xdo1TJ+gBWoYjjgcA8Vyx/wPKxj0PsMVU+9732AwP3yuZG6H5EQhFew
DDIS3+PXbeZYpGbx+Irg1njSY1fpqiHvnscxsdGGCKZvgljU3DYhRBUgaIS0
0sWOXA5feCRMPSsG9I8Ca1g8zgjlOL5c3VVdR/7eFCyIR8i4c0zp1+MHjwlC
O/p8B1mV0gA1DOZ4PhyBr38rCEklUXie3ZqdNhQC/wIf4ZA4MawsAi4Itx5H
wMsIgEVhs8HUbthEVhEq2mrmq94ndqopt2wqvayja7dJ7Tfeqas2IjSjFesq
MOiJRT15+xyugMnl/sT5kf721aKND/diEnO4Qdu46df8Y6lqynXuf5hXO768
mNPYnMUYvdd/FLaiEWT1R3hxKcGCv8mt6rZCdQ2ZJavle8WYvjghxUA1G/to
YOh276beoGsR6pSWn6EsYTWxtoDUHkfJMeuWTpOgBnVDmHYf1nsqHXELcWtq
ZlQ4LyO3Lyqop+gaAcPRgejCKJDVnxTx4P/wMhj5tIh6pH0OSW8LBpAOb53G
GN5Ob6AN/k+EtBA3d3FbwrEsQavwXh/DuYLhzFnFqZQ7sRDReyBnApJV45ws
4gUB1Rq94qASNuiz67VcLtM+1ZRvt+dRGlMNzgZOogn2phe4rm3ktj/4LjyQ
jBD1bOSrbusxCr7zyPJ1zssCvudo7v47fP74StAlPS1Xvv718feAwCIpwYQr
lOqWu5PUXxMU7UjbHA/Westp/YTSMBtvOjDOiHNQn4ziKDrggSr3+tXZtVBR
04Qys8kLcLU9VzwSPr4l8j7hN1SEhRB1tpqf5grTKIj/feBK+5qUNEZx0vBS
IUfjxuEaaLDj5wHBOWxthTvYVObtbhN6E+W0F9gvKerNIh+/4ZfMANnQT/a2
FqIPlhsIn4+DSeuLzqR4jx52MJ10IGdzEF9v9QUI0A/B0V6sf5X1oIfyejkn
+TTT6OYPbBYRYtteFio/3VaWKO2h5K0m8r2c7lYvfRHv43Fc/l01ZGJSrTua
E1mWRztbJCAuX/yob5k90r1QWHMDyX0lurOG0/6Ts1yHfwGdwlGsX5LBLULs
0h7B6XZEWj3MrDOiq7uS4+oXW64TAAu+Y27pPGFv5vxubxdvC3A1sWluePDW
F/bW1v90s1nsqEwZFZk/Y0CVApSxHbRVJeQYxiitGXEfW5g9OMwzdFtwPJiO
ap3gBffSoyfL7Rop7UQtju/V8kc9LhpptNcyrVvubwlsR/6QlKiQZWrH4XVO
Q/2DjnPMusNawI6Rg6QMTXkR2Ykhx2AXtsNKNWyDczVP2r+Q/SY3ETEuSE5U
sezGLV3sikzxSJ/32q/agobgCpY4IOw01dxJY5FZ7t+CQDT+u/N3UK3hNDhB
kMmqualnVSmVhwBCFTJyd0Ufnj6SrlaqivONJoBpzQaBxxBQueYDr2AMFi3P
bJ3f1VKMQsVYX60dFl2wWp8KsiFk738dHqiOpaZsJp7zNz4j3AE4mzU/PoGl
bVnas0TfGTJ/QHd4yH5vbsosJ9GrBk2v1CUkZfDFiPFnlnLHao0c7c1fDpUv
4wZ64b9FQcWCY6ucVJFvwAATYj8gIm14CD5zEb8V/Gs0b0fr467C4jwvqW+q
S8ZlnS+xo9YuazedYRyh9IVKF1AOWKZaDYCqw+yDjG3tA4kCTCFf6aeb9jeW
upCKojzGOQbPr6pNuskOGBeNQc5jDV6OczDmbnz78rWJlbHunrbQgplk7Ngu
S9QpB+CAqloKGIGQfXpmHbCmIQCbaIgLXGxA6kLeec63m3Mdi8XAzlTX5jfT
5C+Hnbjq25eSwfvaF8b7hxFVzbTMkq2FbaYCQRRCC0IRC/CpeLhTCdMStFh2
VYifK9I5FWY9AfzBVxXrS2UvBVy9pCwtXBuKePQSEuz09wAwPa5KtpdKRIfE
doAkhqMGrCAreQVfVEN+uYBiM7KziSH8D+1MkU+5GKXsrtUkvAsQzT8C3EBO
sIlmK7Q5KzUTsiTJ56K5A42Y1TfXwRPSkmquHAKwczGyD/fAzr7Fa2FG3oLH
ihEz2iKjri/YOV2PWutpCYhiCLhrj8GbEK/3ejK8mc6eCEkQkE2vHDV7XSjv
8XbsF4rx0MgE5rpF5GolzCCQrDpBvzumx11Iw35Y5wiS0Nk4pmuLne2v6lbi
xCtEGG9LlQRSA95AnYum1C8ukcmMT7WIjfsNy91qk1Uy4XwyJrlP2Et2+gTV
+fBwozm8+WGX/6d2NkmGjDHEAW3AtUgIb7cv8jlbfIiztj0G9MIsn421nFay
HITo9QLlHPQhxWR1oXAkbdAdkDeDJ1mV7ARvtbOc+VeO4L9+7gzue3hUeQtP
b4YpdOStZmGffRhcA/6pdu0OUB1/ZlXe/PTF3oKY/+uQz6k7Ltq/EWS6mpit
aIFuSkkFFEtf/hrOK+Y3uVleGAfq808UI4DrE7gxEllepW7yOrYSbfup59En
KXnSS1hfhAiW1vQluOhMThXDc1Edl63uE6vnwANBotG5C4oBsPRowFVD+M1G
Zt5EGMweZtIWlGvvMvclWrZwXuc4Vs4v81HJYPYxIF1C2X2dQba+6oE676Va
8oTSPc63/HQ3rBhj3L+uvix8S7vzGjFAcjnHiLOIY/I2cW6WHbZ9qLs3i9d1
cBjOnHVkh5PVhAP8EPepcoIfsnPzZwXO8aDDVwUAlyst2qT8YX3nrv9qEZwK
S8lbmel087+Z3fYG18QBkbZj8aEnsuej1ZJbgB/oqTxJfIGfYcjmhSj4NVF6
aK0WDA6bTYSAxB668S9kab2PJM2e8JAIj4/LfRjXrRtvwl4ZW4EkThtS7ZLZ
O0zCuZQWTLr9EssXJ5KFFQvZ27TizF6HKHUR6L4UEiEOjIgT78FKAEU+npot
O6alQFZKXfvSMLe1O2C/Lv0vozv+17Pm46HVfBbkeSrzV47viokdgShoReHq
Egnb8KTv60sqguJPpd4KywmGxPNXVUiI/AmuaOD/suRP6TKqCdPpF3R/rEVD
io6OY3riXDwIy/c2r4ZUP55IMWobSEm2NvyACPxJW79JbaNX25EDj8E6rnwB
XpWXEzpKPG7W8/QqXzZsIZZRi/pBs98V6gZNzQvtvTt/xgw2iRmhnxj2cpoa
LpCegLGO+mbdCEb9plMoNjmsJ03ij3Cd+FctjOwFn61O9HhV/hZkQ7DhszUd
aCdDLj2atZzxEx4LW+g+upAVcvES9cJbu2o3PRkXIaKcysYTaqGMX1qMvJgA
4YGkr7nF7zMDwK+MxA0W36e+GfqscMD+SRAEXMp+gZ1R944mvyKhE6S357IY
y7mcp4RogbuKF3QnzxX6KkSmefbdYDjqP06VojRBlN0fgSS8PWDNHpe/7+bo
rgdmaH2ltjnUvg4/ag6hSxlXps5LoI1VyiqUQbfydXbXroMaxjlFvZhh5Hor
+WZI7jUESJrR2cSxlPwIdX2FLW43jDpb/dDKquL18MuPLPJSRoYC8JPlEIBi
IBPUYP/ix430DG1iw9fUdTVOvJGQ82tg74ouZ8Wt8Y43jC7AQVjs/0yLppkm
4ouCPzicf+IsccHyWyG/WrQWiHDiAOFzU1ferGrTxAOaMf8V3qmKe2zSdcSb
Zz2foGCS30rR8+xbPMnl6pRqUfjai4uPEfciQWXoNEB5T5iZdWIsmJ0UZsyD
XUvpjy4PXz1M8jXw8kEdzCkop3MQsumbXVeQ2SE3ZSIZBF7LcWfhgfa0f7S7
jlBJfFBv9ApjAgAooWyVRIVEGc93BWr4XvYPbF+IaInkKkG3GeES/prE+85D
+O1shcyD7B3hAZesEetTHauLLW5adxmQccsmTacZ5xbGApkjgSwIVAn4Tt1e
J3rYuYty97vWOAgC/X1jpibXgPJJ7nd+JiwvpCCLe9CCt++/ayIs0CYCf/eY
cHmasToOSOmaInSKnmNaOWhfb009a0Wc21tesu2lkiNcUULzUn8QwB/vGLC4
89sLide+pDAfTKNiJ2XWPgK5QQxqZMjr79iHxZJouEdh+AK8JwaIXoKHGez4
ZdyxopcNcSIIA7YL3bR/NOS6ZhjHX7yfMICG8eMpnibXPvRNLXJG6SAicQcA
5m/1QALsojjKwqgpcUjCN4V2oVdvmBNuCrJ0eqF65DR/7KDQZmjNUV7M+2Es
oKOmd9LTh2NgZStBBRPFZGHLnaEUMz08oRMdz5sCRoIQzNVz5UxXhYva8med
5aStZ0cCd/gK3jMCfkqNWR36rDq0WLTbdWGYV0zm4uJO2QUAR3LnsfnBTOno
IHsuE4dzj0376xgdVmVn2atxyn8XbVL04QGN/0zdpl8kKIlg4tlH6Iz+kHMy
+pMN2ufEG5NrxK0ROLSp2BR05w5NRBuRTlcL6YAl+QqY6vxgP2VytDMgezB+
t0y73txR9v2x09KDfEExbB7nTV7AvXd+PodYWrvAIZnT/rX1ZHG7S7DbpAUl
jaMtnBZ0+Hnt5Xoo0pGMqrM/zMYbG2eRTCiNnL6DXgrga43wXF11aeBVLI7q
uTFPl7aX1Vbf1HQHoIwDKKOPZ6Hg/yzoGFQNCV35/l8gIaEP8N0tIHLN9Ud/
jdxwU/GsgoFKJ4w32fEgGgyyYC2QOJzXyPhMO8BcoLurKMZCm4GFtCxiH2no
87wJTGD7XQI7KutlO6Th0rcIox8SuxZC9qHLOOOylBcuByAm5x7V2Cm67RZt
OWy+/72K4vj2IHpFWZSXce4FBtDsrOtG/JQf6OFkME3/2F95LMaca7zxGvRz
KZpHIuNyYo47IDyJBNw6efOfd+dqJPA3CRsRfoiyl0SBPDJcn43j/5m44cpe
QYxB61PLuRFDPVQ9QTV3eMRlRTEz0scZw31A2xi8G8PL//sa4WVhFqsM7Jc8
VdFy4Brmp83hsxSWbVkfw1AsyqxVCftsaztopK1arCLpnByM9TwZJRfhMjLp
HFuOpew0vEP6syw0eX7sY4vl9LARPLY9ZLNx9tQgNshLprZykjTLJHpB1gFV
aL3pddiiwdv6a4oKBOaG6eyP8zQpTsBhEs7NlP3AIMwSphio6yeTR9h8/A0N
Mvv/T1VWrnrJlYQlwQ3Qu6xduu/winRE9d8IP7uiwGYIVU1nDLlSAIqpWOMg
vHU+rHEzsBORfRQb+Rit3DfFbEhr9PrRqnfbDPJ/J1iqsXlsqBCkLVW9/ma/
bBJu2YzPZjUswsVsCiGsjj6rn9mXxKQ8zzxvxvDxLW3vTsALedWz5LLzVsBl
qzA4V9b+wbe/mkY06vP3zvlkhBnLmt1h6vWRj295HYI7WGyFFhjr83aXUkfo
zwv7ba/0fFcNWt5NbDONA9x0FfYGAyOCFDeACU5Hc+VP6/gpL4cw1UyrerZw
QyK2rtUgsg8/vIPJT9C8G6vhc4YJAnVz/6T6UnIDXSAOUxrGR+faiw23TZWf
GWf0zH+qlyjathQxpeymv3xslxNWpXtTRcxtnw6uWYOUi1CuXW9p+RZROJZo
mDJf7XBBYvmcxL7rZzAXLam6Rd10W0nxLsGDax7bn2uN0bppD7muIc6g9QGU
9LNmC9dGQIs8wvmeT9asos94AnA0VgoF5im2Nk+ahsgqQkPIJT+4suf58TjI
OS7hBOxg5mO+ojIFgQi+yEK6mAs8nCxEYdNPCyAe47prYhr+I11ptz00HOzz
V5ezDsNxofKtXAz7V8VUUdoQmRPnMn1TEnnAzTb8/Yj3bK23icnT+XsKfWqu
a7u2pjTo2x7gQx6F0wfD/SGfdgKDFl6cHinEMwhiOyXZkrG88Kk+/rxhuBCl
8r/Sfyaquazp45z8Brt4AcBQ28V26hTcbcwl0YkDAdzZbzNxL3tbsJcd2oP0
J1HxUINVJZfv1UbNyH/jl7xA/pZtON1q5/WL2Ql7cBzPoPmHSp/kJF9OTzkL
ZRguzig0zIt/D4FQtB/eqDuRWvkeyi9EXWSHSDbwmNaryyVz4XXYrXNi/rtW
r0rhLAlPoYNexkAWca98atovYDsTriT6d2EtWqoUINjlipjHUD8dAw3Dnw80
iWq/kREAIrBWKFr5oVUOQKnZbYQH8lsmHNZjR7dp0/Oww510/BOLnv4VoUmC
CpN0l7yy42Vlzd2fpMmni2q7cX7fKCVweU27u33zZyIZBCHUWaZfi8C1kPcY
gB72HFDTFciytL4cPtlFtkcNmZubmfAZYJRtPT1toL8FDE41U54hvedNCFJh
M7rad5o7HqrITBiVDXu1wx8oGJIFBw+o9Y11vSYgsoXIiCKCGPlBGgNMni16
+16KYBqe3xDdWmWb2O03R4d03FP0oxyEsjb0gVAI4tx4P8TaFTAXGB1yDs+z
iIxBil2YBd5AoQiOF31WPyIyBxHKPXFjuFccXRxr2uUOzPUnVUuKrGWGO/ZH
iBQfEzbcT4yI7I9zAQLKfb/1XdC8M8qu/DNHoUfYUX6JN5UlAsBoZppAN5fv
9asiq+JnPJfpyt8b5GlhUVGsDGjf3Q1uuPqRPANuhAf/q+uMQT9IVsZyj6Pk
Viy5FyIa+2GweUSfPk5cAfdNYNMUJ8/RKVk0zm8IEOiK3Ab6gNdmFvgv9iRm
ZOxqdwJsRMeMilLNkJ+3pupBSiLoeSORkuJCVis05XwqQ4fzTXCs5/Dbm65e
JGKH3Wguxq6HXs+W33NgM8XggAgkFHFpgzl7XPOV82EAb3gIk8cmIVDvrBkh
kqQp6W68sks6gqy9i6R9cVEQHvCE8JytUIowiik0H4xYZCnQB4NjzgwwpRvG
UsD1Nrzpyx8mfAPLiQVF7ZmkRhiLtzKqKTdAQADC/mI+hy0B0BIV4Nh6tMIi
WU8rdsmrY27YrtQz9bh7g0Tok4ZUpA+sz8+5xbVsfYnEt1lqtH83gDwGHOrj
crpzxBvMow0P24f3xhAVRbLHzfNnWMdV3RQ7ngX52yjt3kBO2xZefdg7iqHP
pdpl88RIqAaMy/yjnOCfn9Sk6uci7HA2NmeqmNV0QFnYxoVb8DNPknyXtqiD
QB+NCnTc0DDFhSKm6+YfriSBNR8UY4nqqq20iexlH0K+xd4cVETlqU7rzbRd
OXVzYNhiTPyrb61Cv/1p4EhyfvOgAhN8WJ997YLwMUxs6PsiIO46PtL86fB0
xwzPtqNelKgAyHiP9/D2F7HeYCy7uqf0yVTKE9czCweEdAvSC239IMlpS7ZF
DqhB8og25BJYRIK0Gdewtvt7ejW8R8bxm+xgLD8JPVUlpuLel7lochujpjXe
e90HbAO29tCGrYWme/MJNQ6HcYhRbTQBCeGfcmCG3JOU2PEpdaLs4ddonuwJ
hkecDnrEpUaGhSxTed2qpKNZQYArgnV1yt8uWtM2M7QK1fgrxNjPy5RV/vg9
D9cBQwE29jfjM9N+LsTnUZmLGV6gKpCmDxFLJQtvibnK7WM3FcBY0F1AqCfe
SszpC0juLEo/QSFxuC3qDhICJIvOFAFIW+PnJnlrRDQilOXcIRtuivABQoJC
Med465ArbjsYbpD3i+ZZwFKLqC12GNIxDEIOX2BpciVBQNoqLihC6dEsqYQ4
S9qydE/lv95bzi1aSUZ/fpVdMpfWI0GUpzn5zhqW/61QbT0ZORl9+oR/doiJ
axiQr8aUteD/7dj5L8Zddx9BW7FE82KZ6t5qhasunxKXfn+ER7qVpN9dCCUx
bCYeA/aHYEbQsgL5ENXbG7JhiF3X2p6xweoByYTamNuqkXlflVOTUUhQcaRb
vCwzzKoH+Zif9TggyrSeWL+P3C1qdewE6Mmn2R2iyNEx3H3arHItPHObSY3i
VgeLWTifp/+nk32C6N8r1KzMCAAoP2UdJqT7c3dSAQ6YJQClg0a7d4dSI+3D
rwa9mgUF6Oqv0CnmPZGMHBAiPoFv/FETjnI5DdiFR0k3vk9ca+Zfb6jbhq+z
IFa6KP+vZKaWoGkYf1L9FFwt6bnm/ozVXg5vw7Qo74Yhp1X4ZNefJGmEwk06
Cwb9zeEQMh9VMXBhlzIzG3NHMoSGtzyE6N5Yon7Sfz84HqvUXeP+iYHgf+tb
8k7HdboOrFmbgIpNsCSGyTemPeCSBN6uT/xA4LwWdxGC4z20tkIeW0bUzquF
BiTlySLsj81G6WchrVS82BOxFy9uvWc9WBoDHcTEAo9ymMlvxCB2tTVhA0SZ
ijM6heuD4yQcZKyLzfTDtU8KQv3g8jO9EWGoNP5wlV4hPONwDMUfph+2oSG8
Waf2LZTw3cAr3Iry7uDcqa0e0Kv3aD6cb/pQewTQnGxqnbWfAvufTI1AB5i0
zsrVfMBhFd+IYzCdlQPA0iwTH+P4LiA5EGcrpo9kyBco8RibylHpRRe+GGXa
8R9ohqOXhzHvQGXKfOQMMqeqOoMiqIlYcBD5RNTIVquBdpI5g/eNQFM3/6RE
I+wFSFhOQMb9Qy1jjbq9th8jxfsLYAxUk7Ap+RuEsN2x7QxWqtyDkN4M1voH
T/E3oRHKH0k8T5xj+P1Txl/+1xGYqwmwLIj6DtynJidVE5xgIeGh9BsVFiVx
E/YdwCNRSaYr+49wc7NUOq9SKWrHPgWCReFW42YwXtvqAyXs0CgoAjYdD/lv
CBeE+vAYLSbkak7QejCLEvM6/1vwFf1FkCnK3ddW9ZUFM8Ks2ipn1acLGgyl
kobqrwd9gVywJ6mBIrRs+lvHO1no+4U+UY0ZG4wjhJtv9QeDBkJmMESQGF6u
BmxEM6GxeLuiKGiAoWgkXEwksvTCdSN+HrADOk0Ua3W7Ufay606lttQKAKdt
2tY051KxTAgVnTYx3WphXdiMKPdmbf6bRS0JbEfvcXTficx/RIMwDa3DdSOg
ExsZY8vMb8VTue2Bb9zsjIP7MwSoqqUlYD6N9gdo8qXtBT5cWNE1wVgymgfS
dVc9bUjeaQmHfshWkU0AJIoHrNrnJ/ygsA5EAt1o6zTo35/P+8zqD17nLVSz
VWMydPsWIRd8ifapAE2PVAG5KujCHjTVwHHe3mLIZxQJ98h9NfC9aPOLkCc7
gOTTGR6pVu4b2G6mQSPupuXoBlJLgHEh6WfvjL0VVsRmXC2csmiS/EAnj8jp
0vCRWWY7gpZsG+IEShDW+wQMws2HRfkkXdEOwSGetSm3ToVNwmlTqFswbABg
O1+cPRVjj6kA0pqGXVvGoaspa+SC/d9fkWNj1AQ15fvcasqsmap3nXDMMUHw
deS92L/O0GknWkIr6Op87x7w0BMnCBtz4TkxIe1NV593fJ89vUYdUktB3xXU
BbPvLXCY0D6/mrWvRS8I3W8mz7dIEemAGnhygEgyZuIjM/mc2qvu4ymgxOZR
lH82V8/mgKBKBzLwO7035SZOce6iJCB/NcpxzI1eA9s+rUCvLssO9p3jqL40
JluXU2k6klk+C7k9ZVsuD3rjPCaN6U9k7eKIzreRxz0gPzBxGob3R0sXMVo3
vRwqAVwOu1PuxS5ScD4pxTnNw2/ktnDNmk5CIWLzEMeo+/z7AUfJDBnGnVWL
IGkhBBp4Ds9/rz75QpMiK71tw/PcDBNBxxJ/AdKvZ/mDnfNDD7toZ8Fldb2w
vq7myJ2qDMXB9vLt/VkYwt9lQxIJw/NGKJDyQWB0F4vnWnvHf5QUFdfNtKQJ
UpAkJwd5VfRkUt9l755fy/EwQpki/T5jMwp+E04d8yYdu3OUPsq8nKk4xc5p
jVLToCbASDnXZ5sW7TD72hpBDiUbwV3FcDNIl5O6yFw6X5RVZpIaSxGdZkYB
B7M5C/dYe7a+6EqXaTk26VmSH2lx4/9gY8gXOID/VsKm1QoMoCcwLYUjY0Ul
VLolYN6NBa9iitVnqoFxb9wa0eRKBG5Cb1ixQAeBV7LKoTPwQCvQycaZb7wC
7KxXtUtidPRMvuXZyqev8RYcYKNHLvhZb5k4fQAobgZNhrQbvqFm4EtqZaLJ
zDn3yifWuWZhkZgEr+qnSMpA97REPzjEMok3f/kTUvBbkWZ5OCj2wL4T2dm5
spa5IwVG7jM/jYRl7C+PFhq2nfRHEnYpN3FEWPd4eNbzjVxpSI7zR3qIS2wY
6kko0knBvhSD81zu5Pm42BlRYiREh7K+xdy7P3S0UXA0mK30DU9bKdMitWXD
gditST0ZhUxGUoQ1vC7V+dMSajAs8i2DsdP87c5xj6h9zqfSFdBCKlCC98A2
pX+lf7c4pS7E10OkmQ2llIBRdQaMYJIyizap0L8mZTNAzAweHycBTMjbx5Nb
LIuZahE5qafQ6Z0UMVRjIA2aFnrJcZclEWzsI5cFIb7ztpmZXN70sV/kR4Vm
GBGQcHF3d0FeO3kDOtoeb5Gt4QXYTrVaTgYV0THQuRgIRz/o4zsrGQEQOdql
aUNVNNh+fxMKxPhN1Mi7adFAe0MKO5jphizy21bzmUJ5inhQDkKfc6STef/R
lcQ35RlZsuFe7c5lclPltM/ScMz18JzK4NgSsR6Ap6GVSfnp3E5KEjXh0d13
c9+9RP54T5d/PFxbbYV9u2ku7uz6dd1a5rcav2RRsWPOIBITT1qC29FocVJT
aGC/PF8FuakMxFHCJ3gvLe7oIP6UuSzxZjZDrKjD0Qxz9JcepdRhaxn4jdeU
hPSRC2NUThQ19W+4EIT9BWb1IlyV29hdcSMEBu27OM7lrB2BsURYORazxmDX
EGJu123efpTI+LW/KzkW1n2v5PD1aPu8wN/+jx6nB/7TG2nNzRCYss2vLzYI
JPq8dGWPqDdZVXAEk3UQdutH6FRcBVXIc0sP6PpAd7/7xctb074ogTxVXuAz
08xzi9cdKHOyomTrL2QoLIJuXmUT4jPoUN6K3Wzb4Q22f0Y2q2WyISBDQS66
xGxyNn1FfSTbI9JnMlw2xYYLXssbeOfSMEc9VQl+h5rpJaiR7U4oumJMFGVl
wABeDXWrDbuvN4ugQOoFa9TjwoG8MwMZvpDib9URTyGHzNlFr9xhSqiTlmvm
YgCFEY/9/sZvtQiK8DhIdQSTf/LAj9rD2MDSmX69QIFqseEaiwBA6VxTeSiE
KVNf0nBDgtv5/ThcRM5HUdeDBO9iytFyHxO3E+ZXl/u+PDPqbnQ5mYkiY37p
+mK53h9cvAeHtYfksfxX/VKHVtqF6AlcLXoRNVCD8oS6t9llUjQbSBnfhF6Y
RUd9SYW9wFKvHyWLkUFUaYxK0OoZwDqP0WeQEzmyepENkJA5QWT7811ZaKie
qcWLmE59qcxAn8eiMkU1Jmrh6b35UQHcorynEJcxwFIOPXU4lpcP35k8gK5P
MWK0dxGVV8m7qmeJUk3R05FZ/FaGZTFM4gLLRNojPLFiYYNI3tj0dXnQx8io
OtBmpLg+OteejGdyUL8ekB9jKxKG5XMxbJpEOOQP1WkE7evdjn6ervf1O6se
PhdgsQ3cAChPTgosRCQXw4noJbJ8NqKFV2c0B2gT2ypzjENWruRhXXPsG2Vf
AInX1LCNScu3dIme+Ey14i3bmQr6W1IoZZzNnF1KsRHYqdKoXcOCDM/65trc
cE/MgvOVq+g056ZTAsEs+baPuvjPPqNBdbjFgi42Fh64HOd6k0xropXGEIO3
dF0FNYFKNVHTNc7DIiYts5Ij5lankfUSCKOJlGMGS1gZVV2ochkWWrm6cuL9
Ob6r/sZnewJxHFgbf1l3wAwurNKiqO6I+oN7L6kKHfBZMqJVvwbuUpjmWa9+
pMi3kIJGA/kdmFhsVADXww1MIeyJTYyLF+lrtuJkWcBRZWde+1EXPFm6Q+/d
krwdgBRo6v861xMe/GMfBhf4QdWO12Y4fW26rlGui2aXEGfUR+qDBrXvvLlQ
X3gMsEjuV/hTtuF4TZv7Z05Sn7JER7v6EggB7mJwZLLripmz6WmkbBXi8zNm
eA92yIVwFsNaSSj2USRxtHEAurIjpbBZcSI9ojG1SHfGyxtHskAXFwZ4SUNh
ibWWBynXJFFpfBNUao84om/90kq/8cP5iQLwsZ/H0zT3MVHJ3wwgqpVlR9tW
5hDSKPGdqQwBGc9JzBWOSKCNpbG8zq1uKdp3WOiC5jqOQbx4SinSJtE42erf
NgjXNCQpWh5vKhBMBS9pFMfW1Emdq4aEcMOLODyfjMLhbOLCpREsQ3YgrT0I
qN5BrU2Mv3aJpv375ANPjAry7vB9Z8PaCYs3nJnZuML3SXQHND5SaEMUTQAL
WIygvj8M9yVNLgi5klNHycphj4OshTkUgq0nSqesTaaOvQLGza1zq/J7FwTR
5MfpQbditgrS37zzaJ0y0y1V7B7lD/0a4cWWYc/FydLU5nl3nDaOXx2dPQgx
gHB70xxUruwkWSBQXRIwvezMcsbE/vl5WRGn6/tqxT7AkP11CP1AYX2Ow0UE
THGsqaKIi7NsssVtJq5/PAkLrxRHlLHDdoQx+L0BTXCWiGq/IXPNZABcwrg5
GNgocl+CD5zp06046gAPWDO7opNFgQJHFIzOTD4fi1WFJPiQWBpyYJnaTil0
p8oSg1N0lJSWanTYHl5nt188kiWakP099Q7eFzqBwordGxn61/E6T7XaulPE
cZ6IuXBLluLfDaAOkZbGhX29tch5dcHVBz6Qjh86QDPRQmUF7RSgKrPqtcV9
hfQ4aFUA0PeQaYti2+ZZp6nSwQIAJ8OSGIZoLNtBHzTR6FxRtSmRg7NKVvly
83CIppAHgNMcLI/yh3cxkNS+U9HAHyQiVg8dB/9E3z7fM36HGmOl5aWcx9Qc
9SKOwkmjBoD2Tni7DCD0iZINIwiionfdS1ZylDEd77VG0gje0fY+F8eCiGzB
feRCD05NWqLOsuxe1qphjdAKirZsNylQetn9Tv7YN99dfbhrL31Uhro479HE
HdUMKu27m5puskXYtasbx06ExMfOJdtzCxEMCYwkmfIhJBvAeVctd0Ft8Kfz
ymcmumYAwkmxlsR/jUTJwNxAhKJC3uG//AQNy5bTBkXFYczkso0O4+UIoNSr
ShJ+NSUHg2QN+tXJjRhCudVwlmdNgJ/rLBzCH/ZnEfBM2Ld10UwRjXOHpnQK
M9OLTBeYmEBEXevBmYRbnTdoLIQA7/z85vZ949nhmkEb81ve5cVAKZMukaz+
SUv8CjfviJnnCNY4PiB9mO9uHjvKW53VpPY8Xmv2SX9watXBFKb+X9EaOoXd
AwfV8Vid6y3cLkt4FE1ep6pyY71AZpH1i33WCTbQKvB+0u4CaRKGI3/t+Onw
P1ehSg93BaAl8x8r0VlRpyOqmJsmhdfF9edAFTh2rGudFvaq7THbXSbE4CZa
9NmR0q/4hVyxFz9VVoZJ1qvOXk2dS5iR0pTvrlN9tVBVJmZ0HBLFwzgeBeHm
1aX5ymc/BzQ64VY+zX6q+3rjNBsvA2H8npAltgrK5MFPG3+XjXafKf20QdAD
bBv8pgywhzgVi1k6EC9q9e5CU4Ms3rPJ9aj0VyYlH6rX3y4qXXZJcrInPN7t
/S9g+PSN2AtnhapUCCXffXOppbIlZgIjGjmEK0aRzwUVzyGAJf9By/5UaBsR
d4GQ/Az71kMjKvEbhPWtZbvBpY6XzSmLcu0HhcTZkHDisP3vzPRv9z4P9EmW
u2ZDxVC30KrBpYCGBtYXGviNn/i78z/mKu/blr09VAhuxiaSILFJa6FXb6Mr
vWO1sNECVX/QZFt9pMAvsnwW7m1or1YISpCP/C44vDHB5QCEa/ZzD7fqhDlP
E+zHDtQbKhDE7HMwXws3nx4ihJla5gw6BL/zxbSkyWrOLPcYMCvUnYx1KR7M
AchOQ5C3jcTTirhK5KK5EhAkLq6826vAL4DeTe3FrnPT/koD13YaQU0kF6Ev
xiuCJGGbrkkc/+xaMhGXPH/XTrWs9PIVVOHbAdsEriz1yzn6Y7M32XpaFz33
9v+S0ZiQqSTTY/d3MXK+It4zH3lLTQBJh/1zxvC1StdoLOWv+Zl7evA3iym/
L9f2gBCkoQpBVu1u7DaMhmBLmKMJ0ZSN4RbG7b1ECg+OCaHpUjb3QAY2KhtX
dimwXaPS5o9zl6U89p3xwhkc5zKntih6iA1LV3JwRBjp2DP/Y4Q3cxbbEV5j
0a7FG3/dAUVDco6TifeGCJIC2XpPN/d0rsecygqopNuNxurENEc3J76qcFnc
qGQq03YhArzMDlf4HswqYMUy1ftdr3Wcak6bEuUBXDWp6YgR60XoKbF6+sym
J9MHajhMnijM0e4mNSp/FZEYTiMSYUoDZeo4puXeuZ+xu05ZYkuksFnzTBJF
/pb+Ej7tFOj0kx9K5rBvl81iq5HQAd1yJf2oRmf9g/papzrrpgbAfu/g+438
rKe9TTBAWwgHSv4Jq5tJZPqx0b+fIVXqkxR+YcjvZpBzGBqCVq04lXyldK//
O7PSUioupBwDzXY4vModiEFw9vQAokju8BJilmU08pPRKMcA6MMIaRr2a/vA
+msVdkSKx5JCnVbf1zVUq7rX1duf+PfaCaIpwu+wiaeq3oZIfLXX/3HHcelP
nfHtiTy/8fOA4KooWIZxp45dXrOTfiFMZ7X+lzwflZ/cp/SfjqfOVtYUmy5r
5MMtP2NImWJ4+omijm1Mw9UrXXUwnimT0RX5EZ6NBV4TJ8G9VpaBQ8zq8zdW
6OG7CsxhU2ZwannMfRIqKmeP/ReWPmcry07jXjr1mpSuyeHng83jo2VKdqQE
QB2Xv08uHYbwgEqaa4Vg4bmLdqV5OBYleFxmN3Q/Z9EMSoKDlMfeb+nA6vPD
Xu2Oib4/9mK3oyHan4wfUXHjIRsb4icy30/if+wD8tFdL7jtZ03eJ94VrY1B
hSh/330pTlrwgc9zOMXWsNKr/F7ma4Vq2ZaZxbeatwHzZSHYVyP/qVbNaLrr
JIFnfO4aBldcR93vcSWxVM2IyGlerrhAtU4n+cWYSGC4pmQa0p+1h/KReznf
PAt2myDcoN3pgAbpDLlg1XOIDaxmWTPooJStT8XTOCVg4d1pneaMPeWn41Sh
1UBjKbyxcdIhg/ykmrar9rvEqzVNziUypbijQKgbGQdyj9aECsqCNeQPO/b9
LRQDHSpQ3pEphFK8GksjeAbWSXMnmfgKytq5WrmQUTlN1pONH3Wz7Wdcumne
7cMdYT5LmtTeShcZAib1sqAOcTp1GN1rUaxUmwL515f+p6AYzln0DASDnzOy
O7ym1SQpr/RMZQcxPRtYaOEJJKN4+AZstzg6I4lrV6vk42vOf7jz8L8riiid
2k48E2zIj8oQYTIvmYVT5PU9pTYk8+2mk+4ziC+NFWRGw8yy13Te0g7jdAp+
h7UmFWvhACnm3oN7OOknMCM0eyoHOVxSR+L0RDPygtSM3NHqaa7Gw+IxcmGq
LdlsZlO51pMKPP0jgejoUrWmtUlInOpgD05NALuPL2unpbGWewZ/9Y6Ti2UW
6ZB1nFvKQ0PseXqK6jhmAXAVTsk2rJi9YiwoOclqg0g8iKiohkxl+u2GfgEg
1uwlHhc4WZeqIyp2Qc0xx+65V758b7Wa8TBQmYQCz4ja3gyKCt+yS1RuN3NP
S8vRJSDHxrC7+PTNe2wGyz5PfTmHrHwFe6Qrf42Pj79Kv1KUSE8TbQV5PddQ
KiV+30VssDtWbZdUOIPGhS3QhMrBpXT5kAz0nZxckxEDMu4bGkor8aPRQID9
u2JLRTpinpjkNbLN6Asa8c+BLnIqfkOAbXeV73cxDr4KviYf614KqRu9R5oV
sBlrdqiOwqlry8ucvIOcAWiClhMP06PQa0qcRtMYTQjNBMR1bRPqq8O/2lW2
sffebQ0zy3VlK1qCqJbA9XHBjCMsxa9F5h+cyL68PWtHoxPsZKiOISIziE4p
rzW6LQIqohPPLiFvjAse2jt7kkrZt22PFZRN0qDu2hKBzyIhCU+Kshrz/v7w
W2Vlp9mFqtYLR5aqCv7MhC2jf9jrS8NDm0kqtEQ7DC4G0RzxcypEzoKg+TEr
9IATTqZamxzkwYmZq/rb+ttdcX1qi4GNCCbd8eLMsnS6cgDMXHT02PH+7AAN
kJVNU2s+rtVYX3Kkn88s0Dj+6t7XhB6DeuTwN2RiJnTrriU5YXuiae8FUiNX
yriYEsvZCNieWN/UszI43JpJ4H1LSq4ckMzU6q4unob1sIQISSdouMRfta1P
eug1M2ZOHD+e3VH6cx7ljdKEYXnGVSgR7KIMdAgXBSGu8SuLLgokxfcdbFxB
/lJM2Pt4vPNoDmLAErCnuf8lrJDh6xkZCnocT8M8qTCKB9MICWagqb92PGKy
bSLxNgANOMAlpXrym5WeYIq2y7ddO2RwiOePNJNWMgk2r2D6ayXdrBSnIpY2
pkIOFAMYYVwj/YUgvv1OO2j3f4DmDwxLEDqBg9QPUqge+Ul3WFjHyqrryYQX
6s2mjXC8QSLtVxEIxOLT9RLMkkpjSpoMrmXJvrvCOj/FKRPCXd66/g0UYFny
y59e/gOH0G460bG91ONaawzSHQpaYkQnKkBrj79N4dfaEYGA5SPTZYWqZkuu
FxHrjce0wH20joghHOPnO0BUNjHdVnAWO629FFa6DG8J3pKXJQ5jy+LXa7wB
DvNIrlq5/DMWaykh8/1DrZc/5NRnxKuC4CiPYHRg/xsrtT+U8+pqhRqzK8eo
iHUCypVqg/aXiY+NkWUEcJBP5DkCdWyhp/U1fpeM3wMw8nZaKbJTOQcX+ILj
6aTQOSE7UORTWd+F2bRXS9T8T15bzxQ8fx8o0/kIszCbtcOhuJusLYliXoro
zr+KuiQdRRJK66VPZLzS6AWx0Gjc2xB08LQeUfH5aTlhQZw7/TTCq5l+85Vu
aGrYlKmp7hLLYy1ZeAjaKx3GjfJZwhBrXlCgIxBGSvDnWwMjD4ojMjgPxepG
DF/PK0HFqm9DcWfokZPTdPqbZvt6FJlmaiVb146nEdfztJDdpRd8FHlRmPzH
btFJhtvkNL+8gVadipbcC2ka5rRuTR2OWSaK3Q1NfBO9aF4KosJD7a0lME3M
qYip0Ebja4SpSMKBDxbG0JEhyOBTrPjc+FC/P4EOgsgjM75kazRWp9XMtjmY
iMDTerAJ5caNkz/Y4gYjZOGaWBQ4EXVjEDP7WJ2mZpfVKSva9EWWY7hMKEfs
EVBYKRxe6h2JCAk8h1KCOX4i7qrCvHF8bO6JrGmUuq6Is+cDDUJlf/2sKvB7
ANpDhBkhG9p4FZkEmN8yxtsnXz9eR1Cg5DnmADEsGmodDuYye/pbhVytZrTo
4+bQVLFjoWDm0OvKKIk0N98MBzijGLSPVd9knWWUOL9mY8mQ6ndVKZejRMBU
F68dJ+Rg/lSg/8oLtEhV9Sh53/ll37210naS/nE2ihCdGPEdTZaxBPQeQSCP
seGhpcob77DzrCW84/CqnF+LToQorRF3yiVGfKR/YoLF62DASGtS5Ix3IlRo
69C5UEnPpvzTUZCAY6brQBsJ9XHL3IcicJ5c3leFxLnX+KeGtWbCPNf53Jj3
wuMJHb85Dx1rwy/Hk4SUYRRxSILHk6Mzkjl7voFqVB9JXvwJ2A3WvOR0doyp
rhpljSIP9pY1PjKdpd+YjOc24OgTvJC2Mb9KEmHLfkrrvNwH7K0lpGFJPxIw
+JrndY6BdHPEuEoLFfX2hMOWnM5pL6vj+itb+W2UJTS0mgcie8Gq5APqVsRQ
YiqsLYdRPkA3lYzAKj4FFhNOeLpvaNRySMaUmrU9OQM5+H2Ffr3KoEJvTXjw
UbTNxJxzU7h0O7/cturUkl4m+oKI0KKeiD4qZlsUIzFkAtJzK8ZzKN8gmxvM
kjgtkiut8RBWQE4MmIQghL//xFiTM72sfEeGlW5noVfiZVbgjl6u82HowmBv
VK5hoX+GKrdlmi2uYSqmEnaLaqUB29Nvs6HCm/6s+VHCeCTyYJkgQBz91qzN
3Owuqxhj3xecE6/QzxQ3/TKD1KWfUaZk+/Sam5ZfkmqQ75HwCoN0Cd3mA3Xb
gTywS9UzShps6zL8/JXP/ByiSQ5GWIs7XYRGfRt6NnHgjPIAuBJa3DBDB1O0
WjR63djqZjujqiu7OII7Vfo6UmINt5AJagbc0Xg2LVe0yg/FhUGCzcHmvVnU
S7UGchGAEmw+siHUAND+T0BniHj+OtWo9CTnPEwsIgjul98DQSO4IglGMYCw
Mlzr3vyiYpyCZCQ9QGCr2PokshwsAsA4oyx3NViYxdFldVOTLh82CsEsmfad
JKCRhxzXMSjMpBX7PIy4Z6QYAhqLoKVAJP+ZBEvIPi8/Ae+YtmeMpDUIdbWV
fqnvjtKa+057UlZ020KTWeOhZw/ulhMJxq1STQ4HLo1BCDCVDavTrziZDu4y
ofXMauFNSflzaAJhjjXE55R6dbHHpoQduiowr2YsbS2nsHS7BJQSnlDPgJjn
KM0vt4kG93ZNhqPDfALqYlFvbGQKHe4DQfTnUCH0L5SrTFM5R3uRcThOsC4n
sM1z3HOmxml+CE/qUCh1v9C1xO9XjLGhu7Gvm0qEQ3acPLgviXKmzhkU768D
4puwdCmgSsBcVdS9KC0X5D8n+hgYXx8QynrbWIL33r6LRjsTg79R6OTKPXhc
aB9CB99lG0w5kJLHB62fjMxe2y0Dnky232Rg9PkPV7YjAHsMcHxPVeIWwJ0P
dgdR4UKrP/1h3dJx2wFpyiTEA90FnmJh4ZdaADRsQa6AbhHesNOPWDLnf/KX
zsyB2vylE+wiUSCmeuHnLeR2ZduF+fI2wf1X5OamIM5U7c03OwHuGOh1BVkC
tdT54k8sNH/et/ULRcuHBL+IKzrk149eg3+oXJZoVHUsaOVNGEag+HmOKdwX
v9Z/cVgPLDVXhf7O/RE34mCs8BB7EEHXZbC19QtejlqAySGtactPRXpOEcf7
9vkf8x7fO1/nxFSXbT1jwjn0ZVI7TaUuUIDo7jGrL45p98wE83Rd5mKBe6BV
BMENC8wZAcUPcHHK1d6uIzgbR1YSJfvViAneNdoiHLBhFWT5ZKMXfUHNsJYx
TL8ldl5dnWEEK3JGrjzGp5rV85TgirRgNdAd8cw8ysBX1tvD3e22sDqFkm4q
SbdIQbTl9OeckX9dCHzpKtlGoR7yF38Ql95Zg4J663w2/ICGY3iC9Zv4vYY0
Hb3dkkTR/ThT11Omfqd4yseUQGqDQV++m1Gxm0za61Gitu0VDJVi/CqgQN5r
K3ytQgLsyxXp1jAVfWxdnpLZNQhKmJYn44LdzurxotKEEYgHoFwQGHJqmNzE
vIJsVDHWszPVfLLPcbhcVjEbCn9GvFcSZ2LzdzttPrWLWRKlSo353ugATRLH
MdOSnsXt3Xf7eigg6Vbh61iT8CRnNjzMQvI9giXXfBxFnaFM/flo5hEWXDTZ
1spt2jdk+JkDnoJz0bKVZVxD+Fqv8ZufETniOz8bNR0UqcuMMtPZYSS5LVS4
+iJvJJc/Pw4qQ2K7g35/Fm3ja/nl0TfcpfOWg+QlFfKPOogADuxg9Q1qZzmy
8hI1Yh5yx0aq7lQKiA+jWAUox6eEHcay80cZypYL8PjFAJbIovGlUBABDhTS
JUjfDdgKxGkBC3rX+RCMiLWIeuxKFZ5863aAKScWjz6iXsJ3Bl7wycvWWnu2
mxBhp+DpIypP87GCb/emNRKk6RwKQ1lIeemKi58oJy36WdZClJz5pK6BaGUV
HIom4v22jWR+HoKkCPWEJijSfbbCQ0XjZA0tgZgzaDePiJIPwEaHrS2XOhVZ
CttEN4QXABcWeIHntQSyxtIcJSzK2XKC1s+5Evhnj6M5LlM5LXnUslDwvHF+
E7BFI1q/igVy7GUJBLbIrASbZ3f7mTTNWRdHlZ9vHKkRtwtDLbxgK8maFWm+
aiuwaxPyM3YMnzMiZhk5f1YOnMrOovF8Id8r9/AQrEbTzkEzgj5t/awljj2T
jjfnndxpjk5qTK5ldIU5KAon7x7byPF47FTRWP64o8xfLJR+Rh5rOIQVTevA
ZfthMj/anJeAL2EG6yiIAC19xXpwSe4efNZnNBfDoCAJXTnjEkykqwoIWMDP
qjZl7R721OnEAKcWwP3jVFDhAlvKtaXs1GA3lezgCr+B4g1R0mavmKAfFv2+
WDqoKpxTFVsD2tTB2fa2yILFB2afmoZQuoRkwXMXtzXmgY8XinVr4YmZVTgW
Hg6CygQhHt9nGbBose7wl8bV+dPphuPycIX5095ZMsyGvaIHOAyTOVC17GZp
t8PzxmqGXRByutnU6u0t0j+aR+J0kE2HUA/3JVYyvbCK5jyett51Ro32upkO
4bzwVZ0MOj2OKqEzbNeIdEkNRaeQZiS4IiUiT/RgNJc9T76zI0aH6wJt9Pvs
lLqnerxzvys0h5ne6g4M1xB5FIyBQHWSPO51EEsSxol9uUNnOs3tsjCtuBR+
UHaXdFbNVbM/3rPcZwYU2axKCue1OXDLqAzvnQ95DUViPKCGdTNZYzQougBV
nFI1XbiHJBPiX69Wru0Ge3q4WBcGQrSj/mW0qVJ5dw7LrE/4zFLxoAP4e/Iw
ZHTCppGx+2FNPyloX6xZeb1JQ97JUsAUUDTij9kM9l6O//j7coTxlNcsZt+9
YZxuklE+4wqQ6sAJCc9jdz9x2COgRBpNSjJJV4q+HOHpaLG8kcq92LDdc7HD
BALW2qBbKIxd154UiRB6/GHS0MjeYZxryzC+Xtqrb25xC2z3izXzbSfW5dsQ
dcK/xnIwxFgSFu7UttkbHz+BxSB//Kv+DPeXP8b1bYhIb6hJQPPy9LJwhfFs
oNDKjPe8KZuaAy1bUTWz7kGy11OcANK+mllkIckwo5dLcS+EAYF+7VW5mjTi
q2VzN6i4KnjJPxuwYBvv0Cc0ZOogYf/FmqpdkOaKqjiMsVQnqbR0mHuusNqW
3C+f4optY60IR4c6rx5NbHT2F3dZ1gwTn3atNm4K/DdRyNaPxy2fFrFAE1lT
Rha6uT8R7p9kWWzmuIl+3kNZAXPdZiVGPMadLQYT56urKA7Iw473XPrsT857
ypHFtdob1wnxu9oar2jKEVoca3GrhIIXOf9B0jJ7XqiL+Hjq6l5MUumRh7Si
1HeZZHEyvGDi3jt7Mqn34cZLQf1wMue2vDNWN0FnNLwJ5/+IaLmMtB30vQQQ
afqFa15s+CUL7cSzaeHbmopFBvVhorABvM5jHGcruqKdex0a7/Qmqgx6bUQD
Tq0WaIf2NcdOMRCawAYWaX3nqJurjJliro0MlNfvtVnHabLRp5N9At1bfp07
AzAZZfJTn7qdsxX0Xl2pU+mj9T53ZoP9tGzaRCu5zkV95Q5PcK/Hbwp/gh1H
ChqUbVmD4jdVCKQmlLzeoBOEyBvgb7h9B4GrzdGmnAOkc/AUZlU4ir9pruM4
FCczBUxFA2Yercgcvht6GbjWk5X6RH0GDSi6YOKlQy9yJHU+1shYiPa5u+2L
uwUyfImRqcdSuw9+Js3umtoglJXRkX9df9tJzu3XdBF/ySK16CAX0KJoSRTc
ezB9QfHk3u4Zf161i1eAqH9BbHc+oyWd2yIk/thZ3q6zYdWGGxq623f2mR+J
fCaugqrRHaFruQJgY7RTFmqoJqmvzsWsRERXTDQqhpoJt8AezzyavOlRQwtY
Ep4KSbFhWLyn6EPmZSad3ieEF1/WCwtVc0rogF7HBqf5XrMrt87HsYmIQZBK
Ds/M5QQie25rTOZLtlV86xcUxikksOj7/MBxo5atyoMJOOesAwFgF9xzL4T+
TJuTvNB6vK1zVWIggUe4kGE/RkeOc2w/xsiMWbzuVUlQjCo+jquwoodparMz
hO6Ctf/Xit958ZFiXFMJxq0OsMvYI+08i8KdpnC2tvOSp52RtIrP0Cfbl4JD
IOwQ2fwhMLJVGPSENy7nc3amP1PYq7SVgBwWoAhPxhL1tDSS849VMZqyjOSr
8Cm9ddeEq/WK9ja/7fOaeRioc+oIBA8o5xvIJ47ww1ac0dxg+p3415oh6soh
Zox/UmPRVmL4Qh2ayHJtr1bJ3h2O+4+6LAl//PtG0RHzOA7Z/GQaPMNh4iem
Rs8qBLbuW/2NcMYEIkYHX2si75f9YKheb4H3198aJafKPo2LON6iu1NnGq1Z
8FOz5wqc57T7vSpjh3sPBNy6U7EQlySrJQJPw4NpRJ5wbQfYPgOpq1y/GwvC
MjPBZqNB+nKICNFRWge0nHB3ClfefAQ3fwiwl16Js6qLMS9HrhTqKPPR2Fd7
a5UIJ9MFiVxBgf5T3wDLs0+wsy1H/JfzVeeSa71YZUbkoKNrmeQ0WRyfz3e4
5yt9EPBYiHmeVxbxujojeQrMC3iB9RAtylj/wm9TOgZK42dayyczENvwrSee
BuuZ3mYZrd2nKMEIlXYyE7oLHU9S8xkSHKEa6JssZtjVlr8QarD6jGGwpGti
mmjkmaGXK97NqiKIM69e2dbJXBEkX2VCJEQfQNQQSIH4P2qqXXC/7ovzPNjJ
VZlxvKmQsp6hxAY0iWrpiY+52iq5w1U4CE4D6aXG+3fsSEsa5FAJdWPmHqx6
AmKRuD6y2rUhSaWufjoDlPnhcYaIyaKRh0aoG1tDVaEKFGu9YYWw+X02P2hB
579RB3o4S7HPhMap439eP6WG5aUXSVbxHL5wr3rquNp5GiZc00GutRqW/Nep
K8BprFpZlnKqr5teb7A2OoHH4AFFpT2IQLrD8BNzT3prTRQfx22/nkF9IXhX
IKV5dimkfk4bCeRi59yvA4BZlY2c7p1lq740zCC/n6m2VA6GB0gV8ARKkpmt
R9E9bge5kyGRdsQYWTE9BSuiwP+It8p/s8gLqwW4EUianoZfdaFacLYz9BuW
2gq0lk72sdFZNoVJ4Bvn5oQvcY7oid+jw1vmiY75uD7b/GURxDJXTGfi1exy
ihJdTDEbuQrNMxIuPATAzrZZKTbyq+MuqcPZ+XHOkEWZZHBP/2SOecRQ/F/j
m4BbLWK2KhPvMR3LlrogFDr/4M4Ce5qfWGlfXohvVH8xPMlID8yH7/KFlvkA
UTUaSUNLxprugGrF4UtnsiK26E9J4p4jRw8a1qP36VL0mg786ApHICWkmX1U
aXAUKidq1Y3Hbm4Zgpk0QvQpHwmAYNOwWmWmK0EkI6STCbmrWFroHgWBwUUJ
/QyC0Fs9Zh7T3kW+/CXHzNKk3yoHboqXYg2nYuA5B1gPiq4lRFTC4r76eLCe
83A3YI3porvzvF+j2ju2J4smbmOy8ZhXGc4T0LlJwT3Pgy7VbNUjEGV/17r3
qGgTIKvxPmEpEtyP1NHVdWBjJLeDCKZJbSjhIgi/XPqv5mKRpkflPFRP8Rxr
4wOkgQ/kdL1RYA9l7S2v1OspY20unGWXvm/p1a+Ufqx+akWmMwvwwAO8Qv7b
iaROMDdxTs2VWz5UoeftOwXEdgE+udV7q5ngQZ9PrYC+9WVJdk+22DplU5N2
UcV2YNoTc4RHQTL1gYSnd6eTbcOSDrI/bys6WD9c1fLx8StHDE0xuyFJ6H75
h8p+Kup92ySu+bjodKLE9cMJkBzQe4fXTF0QWAXbDKdAHzYDhcJiunhr1yV9
4i4Q/qRtnLf/UIasv/GhJKGDF+UWLAPyCacPomYZWxAMIaX4bALS5FAaIq04
yBXBIBJaZTQ3+i1zhDF9HsNpALBR5dg8//D30vPbomX8p1het7G+F/rOeufO
a2Ykil6JkdXUXv5JJixpTs1KN882z9wcIiTdrKA9kGl3InVm4A3GOoDAH5nf
5aDCiD93aLGRZC6SfPKJy/RGNtBzVT0CeNjFKkLHadV+KZ8KGLZ/rekb/Sp3
RBrbOST+DLhDEn9AC7gqiM/fuXFAFC+q/xtNgaujtYlsG5mjZauvaDJBorq3
smf7Fgn+QbiBeeV9t1a/aHIvY3HeDokYdGHpahhDuywZ8SRzwYHpnl8ZMU8x
XvWXEsmMovsFwf+8L5hyhSrF/HTrELKSm1kudykulKOzHM1+fv/lrgweI7pb
Rqqqk6wkW2lfbmcRGP+VWfi6NmJkUMPkSXavAEiDpNsHmNoE9+n/GtmHZVyh
zWAX8j0WtAo180Pvcro54Zr0Fl3rQb+gfdsZrkXPqrCrqC8U1CXvFwWq8Ejo
lpHlXDQl6Jv3q/DG8WA3WaQ2H4crXrL0d4QE1yd7lRRHo353R8Hv5DvEO14+
POrjd9wFgCRZrLSYZowh6+iYMFOrfz05/yTG38KSilDZsSVOFB+VgytCssQK
YxUo73ZxZSKzzQ3qPwr5T02y8JOikXWVr0xjrpZqLhSovC0K2+ka6G2ZF2FX
H9l7FXJXaVVT2QPs20xFw20l9OzlGLLQ0iKc4cWjDaT3djuPfN+QOPD3eN9+
//nEAUvI2C9JROxtBdjo9+RmrA8mYI0uK2sjTmLhmi6msUYRrjiowByIsanY
HvCs8sdOe9PaQtMFn4HYgz9BDcDTShmO6A8QZI71gA9AfEXyaf8nvaMXVft4
HuOVdVbBXB97xXlL1O8bHJx1UYrx8rLoVg1g1a3eLLHslqeszIqfh/7mG21A
k0heMLIznVomC2L3BXm/J80kzPD0ydf4Co1GbMaBudR7DvtPR8kzfoudexXD
cAoXqPnPlUY+w+b8BPlcI+6Zk+ryZZTr/l78QghggnByoMNDZ3fMorcM9lYf
gbd2n+8/n+VVadxa+vsqe8UYJbkqAPK7CO7Uv8y5ra9rF3gE839Gt8KU+CU9
HdGBLvvSpY+O05KVslH2UeJjODPq2JAKf067+l6BaFBTqwdbnEEslUrB1kC6
H+ynF5aTrdnPr3Bw2Lj0xf2D707hEBdKAPH0IYh3Jm1q8g/C2UOAjoxjbLmb
WFa/W9UUaLQq1RBVsqncU4e2JOeBrBfoN/mnJzdMMJxOh8b+iyv9ZlcgTOvt
UXonqvzh1Ydtda1Xn0h+q1lgSSADlB8d7nkCbx9UZ/doRr+9yNAHgo9vfM5d
oCZv6FizUbVgmsFNMdP7t26B6Wkft4bU0+6lS0ZFXsO/L2cnitMDP0xJm5LM
Yy7wcq8MwvLltI2joIIqlIZ4XWfCqD7Zq/fmsg3I9Js6czs6w71b5buLc3a+
yWKOwlMtmWf0FCkops9i7ArGqSvdMgVgNWhmaTLmfx0+00vevaYEsfTtZOoy
kUPUBdpdSJ6+zXfXZCRTFLkoQuDZ/Lno0uegVByn8QxX8emWevGKHhgCwKIF
dDR3Hff2vPXYVBo9Q72qN4s7rtg1No+g+82advPSUdO0JFZuA2AEj2KxU+2o
C/KZelcKWD8TAlCwptalv4odMfBn739VzwGwpbxg7+gmTm3D+eybuvMsggs2
fs/uPzbfViTsdSmP85sp9ET3WuQ2dveND7ABjFqizTq1Gi6eDJUIyVW/aRio
wj6hAuX4YD+I/1r/9W/qi5yOwsOuqwCx2I4SvU4nkM29Qm/ciH6tXVon22/M
e5tF33Z3GaCnf7JZMypSRgb1DbpbL0pMnJcUmMzzh69tgbYQTPpiD1fabkZl
nxp3T7bQbHqT1AjHYR/BIrkyxxoVldPmtY00nTluvdxeRMUbRfGco2+ER296
Xy+YFKl6gyQ9TNwvkSoFl2WZIELXRsHxTE8w8XB9R9I3Fvq+GPzZG+pKlekA
YYT20Ec8s1D2EIcraSGB5glnRwmcOdrXL+Jqef3eiDgiRAhNpEKJleSfDhzQ
G+2/oldRl2YPBzJIMon62NsUgzfzT9A+yADzIkGXgTFg5lHpQbbSatj3H4eT
i0NEfa4pWSVXRX4i6PD3U+gpQk4dsbOJCQiingGweQZ0HvkdxNzZY+qbSW2D
8sk+frsmaEpCPaA9Z8r3IsE4r0vl4ailyn/+HPncLY5v51ImgqD5XnRBOcRo
SjNAThhljLIURg1Xyer06hEsWjG0CUBWEJqpVvAVEGQS1Wwc+5peAID2lAjh
btIbRTuXBlGiJBnvUeJhsmnR+mbzT2V6O5ZFg2zNmwKFT76Dsg58zJX819FP
kGWOBv4lelCr7kaCNK/jslxbeusRBvWw+6c1OzhMnG1C0rOUQjCGGQJLw167
1XRjHOAqNxBo1IjUGIxdHdyYxDneNkcu4LZWr/R3qH+8MhLh3jaMTYe/1PaZ
HjYIYyHK1Vwli6YDHba1ZQ70f3MxZxGT3Gcv2rsKcVRrmUKYWZUOS5xXhuxF
llTX5cdsMnrbQrWiUWI1ZjNBlrWztTC4D9nzV10NJX2ynalSRAZ4+4WXAhV/
uc9wPztRcPbxTA9bqcvKSu3+1wEz+DKxatsEJwUbwUOzbQSHmo6/BdeKqfmk
XL+5YTcWE4si8l0YoNjyBVBo1yTHL/zZK4dXMtQ6ZKAEBXwpmE2pJSSVVWSW
NHDIHYk5s3fJE35dfL0fiFKtu5hZQz8TegrFWTQe/DMmpSTG853nSGb2UrV4
bPTMln4HWYnNQ0AaGrQqtHCOLX3D6cA77MI5S94KslMKICO+H+y+9rYh8poj
sonVr9tP14yC7wEk1lnfFiTi4yF7txXFeuHo0RfTq6dVXQoiVrAsNNEkiJOx
NV6UKWT0ymjCbZJaXuEgCAefuDnX1TLmfw1roEDclKW2zfLOWNQW1uv3A9Pv
DF77WAEa65CUi0mx0MNBPF14Z2QSjmwzPsv+cjvpRKd9Z6i/XLhu4/XTgrBA
a9KSKGmylTHu/PpbYZjzPe41niMV0FhFAbrh2x12wKTbprb+Db+fnl+o3Bv4
tmmbO/g/A2AkLdGuselYyLTWFAOfpVpCR8OdScYs5dO2/Fcwgv2cTaJ0WcLX
yYwFdc86GFK61exn+SDx/lvmke3TFkBxG0l0vSCZOtQio08W0usFoKkF4kga
NiU6BH3GOwhzLcUH96wGIY6dU8o83HZKV3eiZJK8mRhQfHtSDbS5qBE+mFsI
+4pjwsgimr/folMSe/mX/c+3+qHK13qWr1I7zCVVlAZTb6b+yxc/iw495fJs
Wh7aSMG7lZZ0IMmfRh31MFs1MKzpgmp+25oDp9w7qIcQR8pclrEmDG/bUFNv
ERnyIx96fyPtQB0UKzvKmd8AZwVkjteQA+sS97kH5K2UBm+Q0ed2i4aAySFi
259FFzaIl198xe+rGH/iUGMTkJ+u+itPjYhBtr5nLclrkDCnkIff8gFHPlpZ
VEuqbcdrdBvKQpju/CRuD2d8YtsBQS7mIlP0EmxnwO2J4VmVNDa1lzSx/yss
+0I3/lLgm+1xsEbHKj4o0N+a3Dst4LOjNwPMP9V+VhkvUD7TI3t7PwH5eATs
ddgop/RVIjQwvejidQzD8loxU/XUW9i1J7QfSDvIxdn9CTgIf89l8CVIPCZ1
7yP5MvHu1b+WzyYy9g3eWaG2wGAIusxmT2VUkm0w58L47uahU4j27ng0w7CB
t9+CDlfNpzK1oliSu7u6zRTCPVE2NZie/HZ7W0sEaCPpM5cyRrWv5D7QWrC/
hTSrO+Kxoo6pHDnK0Idpf8pAw4yeE6nCXIgWlrxyLv2xTVZvHa+zSmK4g4eE
SXetKZVumU1pHmlYsaUlwnB/GD4rzPeeCBcoKdZW56Yts5aGtjlw2w4Pb7jX
vLGU1QWygVWoJQmxb30ABBdtT3QFEpp/V33P5LfshWOwqvu+4oC+4EihapGh
bFIhdLApflr9PTlKIwxNREZfX0HbRZgpym3eWWRh5Tg3TNtSLtySvWAUDaY2
qYWEulBV0a1lZ2HihXVhIC/5glPWqFKBQEHDmoAU8CZnIvJ1UsqYVesbDw5N
1y+v2SI58lKxrWz3rnm662OdQ1jMnqIYGCEqBz4VXN5XWpctA6jJdwjnKNuZ
14x2hbRVJnzkpawdAsynDIhLnGki+MrH1dVHGzHJI4Eb3dPNSJrnGmfFK1Wm
QdcQPSJV6d7wVrZx6cH8nKGc3nkkQkkpNbsl5w+v54SCx//C8F+dKQMbFO+5
WtE+XMEoBiqzfECARJgaU7KzHIOe9dg1NXY0EkzNC2Hw31ZB8Y/hgIldQGA7
QtDJ+YtRYONrqlA/CQ8nBsSyTT05NLTgXA8eHlrW4DY1I5hNuPXDY114UNIV
Whj6Y41IghIk6CARzwbc4UCPrY5g6l1THSzMIpJQh2pKa1rWTsn7zSvvfBv0
KnOH3F+35wQe3a4Bt+6BL/U//yCSdIQ1+cpetTiG1107wGJqvAfAj95mxNnJ
vz8gcqATFqYLe8noJuRdlIFA99sIUTBDmVQWsrNuAef8R6RI6RewdIdB9Wi0
5tKxXT/AYUXWlI4tIJzPfQN09+pJInpQXnFwDTdjan4yt+t4rfKn8HTyjknA
rOiadCx+75pTcHqMFdMlvAdhrgr8sHwMqPZyExBnLkOownl/6B7VH+91qzNE
duJdnxqXmRZOBpgC+OrQ57w0q1GsIx/jUqSoaaJaSLYhaAJ/J02dqlcwWHu6
/jb1MPoGSXdo8mIlndlHWTl9VoGSuk76TIImb36cGisMc68bPe5DnNAEccgg
+QvZYu75CBU7B3KMl0v0n7vEd6Xajc4/hy9/q4fyrKqxzEapYzLrLCZHeTUc
cog70QbLzNgqf5lY/aWVzWgkdCksIPRQGcyAliPy6moXEINE4m1H0ujNTATC
z5vtTHmJJYuL5IVCDTSeHvWEgUzt/6b/XkjHvTyFQ+2iPjC3h9RCtA05Wq9M
byxZXycHlRQkgRNZsDJLPWJEYdwYiCcjPlUebyWWqLrQwQmzO1hPMPLKcEjU
CgXOPRq/zdF8iT49FZzMbTj/gNw5xSjITo2Nrtn3cd2nJTr4EEDkjOTDeXZi
4J6GzM6xOlVxuiYEObZVeIjYzsp3JGaMxB7Q/OVfhYqgAjYcdPX1OFGQkEBQ
IpqrTXW9pkkwaQ3VCgtXrydGhJju6Rp+2Qq0HU1hyPmqDmF5Qc41OzjyrIhy
QUeIVEgY9NHdantfut6GNwRteZRy7bnch3YPIEkzSode9T29w3UqStbJDyxO
Si2S6VlOel3RoIimaC39IE1Xmr3mIgc3uns7Xam1+V1cPAvnqgN0RtMFPTqd
eN1QY4+hgFxqgZZ56AJvqaNaGimgcUQKKn20BwXVpG+muyfbK7trS0OupE9/
HZos1dXnXj+njgF9thrzhkUrq6WYSGzb6lUVfugWMaVLpsWTc30wzv1KFPB2
3Mie/auZ8t/MNhOAG4uH1oq3NqcWgx0RnWo/nTlArNL9E0b/a07Dv6VS+zrn
Tcgoc50ly7KPZQF64yfB1IQlKFFaDsFlbDkTZjp4BS54SYDVvxmJyap1CIfd
ItLJms0GEQAU4QH1oRKwOHs+K1jWsyX8O7EPIz+WKuDdHKM/lQUyRTiTrNjH
kArDTbiZrGijRVFKS3sZJ1TTzwHXKnL/9oDxe8AUlHMbsegnddq390VqbHrA
Jp4PXSCnjsaZ7/dEYhU+ibYY3YuRFk8/Pa8UfnV3NzAmSozOF3hpB3zDd4hq
gFESJKbJ1rLDyiZ1guTTg+JDtcbe9Z5a/zKX4sqYPUJ4PRSkyOWF0WuqEiB0
AC8n/vJNEwEEKv//07DticbBrhwH01AZMSAolRevsCmnNQfsuosAcBoX/uNY
vsSDARaXIUoA2/Z2sh8wPl/IdtGIpGhzQQzNYTO+PXVUBPLURaa/rNq2aNiw
DuxIAexyj9dk8RXqsfbS8Oi9bssG6R9IzIM5zdIhSZtIcNtrcuo65DYtscJd
B9c4SvwQutdQ0UmQqOeEkqoHSct7FWTMN6HCQFeCo/WXvnszF5vwpYQLUwbQ
zrIshKE2h9LMJfaxPW7DfYRu3G2GoRUCeE9LTtPv/JVNhXjVaphxaDCLfJ+U
/9F4c/STEaoPJXsNwTNPKvd2UxZIue4vuccUpq/u5U7sHhCna2+jaYuCzX3J
qsN8LJL+c4Kja5rXq7qWghsKjJKqtgo8jqRHRrnbmfKukPsVXArLjcJe2VX0
46r3mDbRuExnB+4UEjJFUPM07AUiwcw0mbiDjwoTFtq+RPblDQ+YmJSgub1I
2+/h9ZZ1Ftoy0zQtnUvQmcKXMAOwCFMl82jzSvIH7KpLs7WBsYlytzXcagyb
V8whBCl/utn20TF7aHF86VTDyFsVAJDr7oelMOcEx25i+VU01VRkcPnz92cI
Lb+hmnNITsbk2UjKwjgqsdA54s7Gon8AdpdNJfhVgm44cjEOo5M7oh8wpsh1
U39T2WAAZjHFc/JEVaDERS21n1UhTZH5kIrfWQ1UQJOW/pqAuaZEZKOmy2n6
AKWLXifqghZuooVXbP+2C8aeKi8NeBP/dKeh50CHnbpywqAH6Hf6WzcBDkNl
17n50NcEl3fDI/8PmR7x7Org1taspghZ0VM8q/R62HukBbd2EnIkRo17NHHF
D8GjaTrbaOrkL3O5AhI2j9Taqn/4q0T1uD5tAkkxuL9JHZV0bqWuAaS0HAzU
VHqT3fqGG28uK52whu8BS7rrpu9XbMDoOWclCz+G5Kng3D0ytWr5oRucuXak
n4MJsUsUcq316ujhqLpDTYjrr01l5QPmcNAULx+ukkqBVWwZO4e5c6sOdcy5
VCzezfKr1kbpMivGezzVP9o3YHQpyG2STtIGdLwgMvgzeK+z9daX4RxGo12n
gZhloQlLrfp3Y0V9h2qb26vGMCBz1FhN3yS580Cr4p8TMme2tT7Em3RxjSTP
faeZaoDSxN6DGTdLEmoENZBugxDMpXuYKspgF9kzAwkDajm8/CbHbxFTi7bH
F8/YpnEe6xDhAEoMzaXfyF9lKLRSgLQkdgzXeALzp6UaUkYojxS7tBpNRqJh
4iRZnMCgUVRx5UohYEdcgizxqggGeuhlFRYm1fOBqmtZto48ARV5ITZcln1h
CPtpzECzGQhrYzBNzlReeLXwoLD5pTCe7eHbijeTlF4yTrgco7Lx2bTh3pII
bgN5oIMt2evmmMMSjTM4iGXgQDSNhq43jsvIGXcn5GlxttRuSsLPdPnxXKzc
ADU+zTz1rUNzYbAz2iou78bXh9daPsPPRMItg5tINJdXZ6RCa3OOv7huBC7L
9onJkab/DKgu00VXrIaLQovNLyEoengXJX7BpIRpAE6Zaz9ePuJoPyVflMU7
9vSJJGnhsUIHWMhpvajyGk89foKYi+5KcJtTAeHm5jisHMjtM3Z2V3IbPiyN
HwOrYM+Bej0iactCF9Pk5DceDqzFyYkCe6cRcOenWGoizvSMnqLw4KQ/U2xk
QYdQ0E3iCcEGWqgBIP2nJ5aqkxWDCfzuOUbv+0vEznP0Fri69ThIuwRWnrt4
lMDgRNTe2x82eiv1FhO+L60wiMRbcFGQ5KHXCm1AJowuWO+NVg8X9vWH1mqn
+/X/QxOyCHpr21YqZVgZMqftKBawZJXVaOkIKWeVcFqMV3cK0PSIKR/Mrrmc
hCQdx41aYO/h/hsJfIZMzJKSR//iGUEc1TgVGQxdZxsE23AwbLVUWC2e9rNj
MC53SaK+Qp9Llsyi6dVPDstE4s7EYRL+Na1QLR1AGCBO5f1ibrTyp3jWq3cJ
uB8KubOq/3605x0xSlKvGoY8XujhmJeUQFZY21g/DfyW1ijqkB5Lo/PRzHF7
kK8PDyuZxdQALVEKLw14yWl/ZBQX7gSNuGNcOQbPPikAv3QBHX+NjoLAloyX
jReGGSd97br65FnTO02Ni000vbNHPc5dy1ED/rrgMXdzlWsYpi7hEsegwvg9
buGBxvfLeoC06C5lkAXtBLK9Yki8TCcSQM2yZqrtMvd9p4UxYmv3SxpjTbhW
sY9K9zuN5vYajdHupbAEL1hkcsRzdeT10HHWYoKrU6sdcsVUhfq/YubTgU98
kogSZ5BzXcTyRpf7S+K4j2FMbC0/BFx7o33EhM1L8GwVjkt3K+0wuH/497Xg
sBiliDOtTYfyQKH051owzMYKg9ioz5+kqFTDtQK66Sgu1kAMGgaQ95ZiBYX3
QM6xLdWnybLGzEiOD/ZDA8WpQemaUtIEhnQ4pFSAZIwgShjHxdmT38fFujzJ
0L4HHY3gXR+aBEmOhs408uMeQSHbukY/s6SqqKXCUrT0xU2AUyuyOh4sozc9
fxNIbTKR1Ny690vFDYQz/HBYePgrxuRJ0o/YQN61+bzvkRckGbEyiXevRffd
D0mD4KTKDv9e1eSfdZVegSvj3r8r2AqTuA8n8x0WBDX/xPNd5d40hvMbR2SK
aJcPwfy/hsn/g1becunKiLfizYKgBO5tiljrNHsYrJaM2FnNWTl1S+8OeTAd
m+Ha7oe1x6wYgmMDd+dPigJ9mhtcl1BSnZy7rk2IGtxHxE8NnHt80b+k+iJJ
w/bIku8zwMwbaPBrsq/anxX34J8P59IU0HizKWesIvOR9BssIy73cv1c+TLz
Pzd1DaKvI7M7Bq4km4VbeRX3Mhd3H1yV4d/lDFdPjaCIKL6xWR/o4zBuSJMA
FfoOWzuV4qDqPJf9fquphXgDtoZESVRlCGPsf+bj/BnKszYxj0Hmt7DsvFse
WuC9wGBCFWelI53dVUP9kWqGuA80gD5EANbhapqx/k8SXEgQpYdPO6PZPFYU
IaoCFmQZZ9Be5tDDD3IFS9tcmOSuHpNH/WOvkSPp1Oncu1g8MdftRb4JL6jA
/FEDBnaVm6lQB1MwlOIQmq5BYoj/siqqd8pY7HtgIJYHXS4IdXQch7N178rI
xT8xh5ZYHll/kO+EcqIvYcI0u59ywEohuPhSv3REmsteopBRlHqVooaugeIs
cEHz2fIob/uWcLhsq4YFIIZZ8+QHgn87iNq1kLBFgUhiv+tYSGz0qPo7jU4O
WIPbwjOnDjM8rrTAVSAjOEqLWjspd3YdHIQDqaNcpd75ZNTe5wg+jx+En/Xu
pOquvWitiDyLgcUaJwj22emMSLzx1yOT3eVFdD3u3uxpVud2PJWJQcx3NoGU
2pZLGDqK7dhHbGNKozAA4GavdqPCf1Ac0VSAaGzP1unPJ4Ysyd0T+gwRzkS3
tm/Bo8Wa9AAHGMqguwgjNR/yLYg5LlmHM1KhDM341ThFwUfljzJfoRF24lhN
r1Evmeef33//tF9P5LJLiCUsdMqeHwYC8Zbzd5BM8Vktf6IVhkHCJB7dYD4u
uy4Rf+yPjluoNtwk0fEmGzoe3U8boS0Z/AO9x5jQf2+CzbUmH1gy6ZK8swC7
8Kt0IKOcQDSvGZGIRnWTfYZ/pexbJvh9ThkmXdsFfRTdPy5q3IVS+O1drg59
wh6G2RjxHi9lp71F1FudnWhQuS6C30UG3KTIZawmp6gyxzAueY7/5cqqqVeE
3f9e8Fw0oa6co8p1t9HlTkLDCs/n0pef9vlhsv6FCro35nuQn4vs0Ccc4Zi9
p1bucXZYSji8ZxZ2adPRB6tHzjI4G2ySkbrWVg+79saaxFy1VjkbSzjU1wFa
BagFWUdqjZQ2plDWYufIIgqV/9YSHmhehvj0jonSMmwhmRp9HBZSXQTKPPNb
iwEwi0fFQOCsSZh90t57lBCGSATnGvhp6rq/a9EPo7X2gfJ3bg6DtZ2roT/q
JszDM130jytrrgJV6ks3rwSM0BvMtc2p8Q1I0PsHsjgIgBV3bVYu9oZwUrzp
da7QS7O0udfLdNh+Hg9vw7K5Eif7IrW7yoUcW935GL7MvM5O/nb9gB6cOOo4
dvNIW0PC7z6zmB/6GCtykmxIdtM4jSikbWvf0F08GRwJTXxxcx2ceDjdKN+H
+CS7P8kKfC1hAYLry+7Dbt127NpcOsFfPyIAmAd6833oawVAD+68nWh/1Dr6
51YJ/bDXVaNeOHK+zja1ce/QhVRUwF+hL/2h5WK1Nt0N9dftYQyOpy1NHjgs
Cjn5frz9kSSq1Uu8E2OM9Otk8qVMCp6MVOJxxzsZmYLRvsVRIUduAmNce9ng
deChbUWXR5AOyJh7lrYVxefkKpIPitxMkSxjLlfolg3MnctOX3uZNHYD/kWe
8OJ6fm4dG5Ies4VwqdsLxoHMN1CxCVURnd2ubVp1fl3RMqGjJEnEKJGO6G0C
5NdwrJEMQp0zpMasEHXlS6CXDYk5aJHl8NFoR3kfdt2BVOuaqT6G9GxQG4bZ
B0PzgLCltDREwzuf3C7dLP21PAbcIA5r8CP4OQKhSB8kA+e45XXpaJY0AC10
Hmx6ugPDLdpK8clyThGdALzh9XhJ8HXVkCklyEpHGq7hwJepfH0vWiyuhWLR
arE4UmKLF4rnll769MEnn3CzIzucxxfjzaA8+5PdVbcXUukOhHNbM4jKmTwj
///taET0Vp52ipP+wNgBhWQSRe3qyuCRA3JRQb8TRh3bxef9+3++f5/GJ7oB
lSvtcSKKZEcWr6ixwJlea1AnECGToWoER5Et/RWW5kkDA3MIC5bhA+m09/Qb
U4MmaSLtAOJ3PqNuahE2LIwAglGzT9E1zejvMGfhElTXevzR68s6woSiYeL6
YZhzbFEWxRv06bYobT24zm5IEsBA027xyC0d519Fyx+s9xyhwIcLk8sfxlo6
lr8YYWOXqK3VtW+pPMCg1Gp33OV/bUwGqPbINo+Y9HiU+sTyY6zMyrP2SuL6
e7V6tH63TB4Ek7QvZWonxVwKmAZhaF8NEZTykVagYnJ4BAC0Xor3Mdh5rSlR
1/tgMdhoEql54nFiRjbVSDDrTQCG3AVc6ZS/45if0wuVHDHETZEqWKGKzMvD
RfTyecZTKM17Jp9+FpQgdwzyiLNHHQTxDke1iQS3wb41k9YGxON8losKX0j4
e5feTakpxjqhVJz45CarheAtKj3C8zbC3l+g7YGMh66gm14bJHVCKjm5Mlg8
jirlRfpgsnFRSYl0O2dOqvxKgbuY8YM2XQV3hdHg4UY9vDGB0FseD5+zFrHq
Dpts1vmt+uugjIhWimWwYB+SwIV6Ei+/xV2i2BPzKQnTTYiz9uEVulu5baJL
KQID5cp3rJrzcDjxV2xewTSEzLh35bAMCO/AffYP5u/S2yubh/re0Ehuwo73
rP5cMjNny+gK1NT68Qd8JAL8ui6ql76xhSRN2ficD/o0eiYO+d4hgJWewgXv
8FQIzZptKAxhivwW2ZOqFgc/21LxhypIOaO8agTvroDOLAyulTZPucUqEUcQ
MNya9MzN1WiomFVeFujGy9kaPbhO0t1ca5UISXjmOHwB4ugyNJrYNrOsEHtU
0KPoNiYqwvUDIXJKPC6goqLUxW6Cog8vQRfSkSeRmxqVZvlSX09m/TJzeQbw
ywFQLNGZeQhEZdjY+gKZckZY0l1LaDyo/Aybnd9wal6ycs2ZaqvyZFBmnhzb
IEQ8g8s+C4Y8jFagmWLpB5ofhQeBKACBSw4ItmW58TjEgTno2TVslchRkqFm
i5Q7/HHSM5LK9a7sp1EeR+5soS4fdTmc091LoiWb0Z7AvS01ufTSbU+Tn/6t
6UXosV7axLzCpQbE0BHnlc6hQ83RSo16VRcXt813e8lkLmPmaZFwrOCrUZJ1
e8Y9fwGZcXOxAuLQk1nixdQYoc5FMe735259JIjRTixBNKMOkhoI/t6jbIVb
iE6lolHpGMks+oqIN/dghC34lXikfJo1NRzWUhilfLgxb4ai2+T69qd7yyJ2
bQP9FOKVItTegW50FI1gexdahjCsdZFVjiuejGSvwUI/qsGpB1bFosdtPdW+
I3q4K2pxAWWgxJ2Az0kN9fk0WG5e4DWZoienl6fSs/qMFyedXuEIgroXQ6Av
7nbLeB/m526vhvmvMo1nGeOJXqm/nJkOvlXZN6XqHIqZWFRoakBREuMlnZ2T
XV62jD1r8hp4hzlVznGDqUYkGspfNJFwsyeJVVJGy0H5QulUZgzfapWaK4Fj
BgH4Ufk1UwHDcGZkNZWT1OmNlZZ+Ra1412v+9sQS0LuEvQM+YO0XpNUlGfvr
IEx7ecNBZiVP+XYr1eNgHj3+IWQ6wDWLAlQDUkpukZ+gVO3yk/dSF1IMLqiF
kDLpxr7rqA/rD8bLltdOMo5WIlHS+tqwHrTySPpaSX2kUJjglfYR3qHPHle5
9ecPadx209nYW/rsdL32KqvDeOhafzGm2cfCTAANijYQI1+RRW1vw2aKWrqd
6hWvq9HyEbqqMgBxEzNLtyno2lCordH2+yLYf92AU+Y5uuGadlrneKazNMPW
+UkYehnibnwfuUuAoZVYNWziAq1SEX84DwMrJW7u4IyldbJn0Q+0oeGsgLWn
sZkw5QDIjkZDT2hogR2VxaP4FqgxorP1uavANfAb1Sul3Mcw1U0fqzudjdoo
GiAoDhGMjlZScdLNgE+uTQPR/Dn0mxBzzh+dzOeCFjzopOK1VvYFQHb584rC
Suhvs7Alj5nWfPct0yyvtgUUf2G+ReONdJ+R6glT5hD0uowrDrY46fP4ty+Q
aSCe+ubgh58XZBcIvzYvlRYHy/NdoEE3wXFlkMrOYt3Gh6QNb3mIwZ+Hg5Yf
49UU9RFL6rnqHtA3d74Kcx0Z5vT+BMtPycWYllRQsv+iqhuGk8qSKv7BuNwW
1ggZLAuKYSvCW+0AAYtyOxBvgqGpPeBKN0JXtIgi8tSK6OBgvUNPOCnsjr79
kFBLsPA261iXhyaS5kFtr08QgWFeI/USgtl/jFMmTlqxx9qYTcF6MZdl3MAE
VgncxNuWGX5sYCw2ifll76tI5hYBctbNJa6o0s2mIlN8tOz6XoU9hflKuIQh
iBqmvs7IEEdV3JqMIHHPw7hkQylLyP+A0JvJkqqrZnLQFTur4vDMUqzrrHnf
R0oL9ufLOoQyxzgUatZwIr2fyMO2036LVnW0jK9AZW3fWh1Talm8bS5tFt//
AbFVx9qspj9OmIdIlITDge43k0Cg0HXSvqtitG9IqvS+q4di9f7a4UiRHvbU
yYeDt0J5dKOKkbaL2q8fViap4TkixgX9Ab6WhPkU77Z3bpKzEkiV2EqoTMKq
oHL64Qizoop/ctwidI0qzJiKJIMG39p7Q2crfYsGqONY6cS9gWKbn7NSzWR3
5/yLgZ4+3ObY2TfaCpWNYXkv5t6UTaMeYrpzGAWampxnmR6UQKHHLWQqBStm
rUxxBHBGdxcCD/7HB9ScHK+5k1HCfrx3TCFjLGNaLDrtsTan11ZuP28AGOqL
C+jqpiml8qepnujwOWgH9Z6oxvY/eHfGAz79nEqy05dJUF+BYifuhT7Ek1m7
ttyRAKAO3qk5RqDnOVWmqy22Cra317LvGeG0SbG6jIeyx6HRDWvXKEaqKA15
VaDe1yXhEthW8lAm7HRMLySvyCAJCVZ+py1jvgoEbs1+FFdDKGgNUoJcavgw
Pgt5pjvodXqPU7rOzU8pAa3fXKTM9dq6RhUosxzAeOKAv6XlUtFAV2k62NR1
4QvIfzIuNskGccqkihQXwCEp5cb0rZ1sFu0VsFpjZMckHSQrIMLojp3Rnl1D
0Qp7v6ivfZlU1bpX65tmQTX8d2aNzdEtgdNuVpB40vztsXoI9O/1i1SIfaNr
U7dJ9sCigrD3B24YUVKEJOjRQcZcEPhxbGt8znnmTm65JRJklM0PBAgLO89X
AXN5YzAJ0ftZH7S35A9e6WUwmw6pbM/stV6DIUrQbIr92sIuFfKGej0DUzr7
bK/4w2j8hGf5rjv1xb4inrVe+OLZlQ/dUq9ykyMkbpHdXZpDp6T6UJvMWko2
OE6JZFdDGwFuyvat6w3mReWjeUAXxCDUlw7/kEMZ9vr1Zb2c8qMUyXK4Rp4R
8jZcnJmbf0yZfiLNGZpeRnPrQ+ZB0pGGEfKa95/LXtZJEhuFUp9dTS5u5Hf4
9JNx7Et9q2jEUXL90Z9EedsgUnzy3g2fDfcKmIbAPat39BweJJJ8ydOwzEm+
KXFlEEm+Qj1oI1K6S61fqea4Ci/Rh/sq+u+doK2r5xvf4kpdo4/Cbu07X7Ek
s6383keBNCgrF4W0yUxYYg9RG3XD9ZLayFp52OP/DMJdjrqFdiTwuB7kWN3k
EaDaqV795MLWOh514HWdkmaBSU+RYMSgJRNgAbJ+FZAtnw6X5w6jWVdbgv5P
v7BYZ4ZuOcl1OiNB53tD1/5EDi5CYk7CiFvvkJwNeGP6JOIs8Na9mPFnzV4l
1OE65fohYVDujC/SAoXYc9bWPlmhCJmEceeNbQYhcUFXcZSDSVlOf86vQgFY
TeXmBKSN1m6GyajXJp9z7LQ2ZMnCVRbHvjAKxqDaMMkWGEwVkEqaSsFpu77q
+ZSZ+qTEI+4SucreLXsXmBY2rPo5VNwb5GznOgukeGvy/c7VvTfYKbVqzf1i
RgkRaGvvRuu9CJM5Se9Nx2rIKV6xFmK5PB83NW+ieJG5HsbUq5tZ4sIfCNkU
yeo5Bri0OBBMTw0iKjOSRrPlGgbGDUpGUXl+82/c396M15QTPlLItULpBVxm
7KekMQyVDfkWcwsN50KEOgUZwqtDQbnO63+oPpJwsvojqpJlloZi4HvxUObh
GnFnTri7JPhRckgyvT4nybpS63u2aDZe/cvDCzlsoVMJqGOdVthjWaEl4+Ch
DdO6MJIUK8vAzJSK2VD9Fqsv8Sqs6W7IGZZA75tBJP8qTgOycVJ93MifvhXW
kVcMLIH6w9h1/x8C1kDpuYfKzvAP9Z4/6UR+5IAy3v/tyGkIKFDK4gGOITtY
efcdaC1415igyW+dqm524mBW6V0SaEwG9uHijEhx5BEyadDk0C4VnazzaV6Z
ruBexzfQrHTpczezXKO8MmbOTIL+kxB2WuDMf+f/MbclUO05EUv5tbNqj54n
Gut/skj2C63KB2SlIig0Rwm1xVXUwHmXwffm+wkkGj7UZE0GMKPeDqZ1QAdF
9ky4kQRzb7GQuFZJs7dtdT7GdZr/2+gtSlhqbbXRWj8Enq5bszct7QfBB+KA
F70lWDtdFuS5fB2KhXKg5j//pAPXMXnDejSDBUFhb5SSW9Wj2O3rAbqX5CD9
WoXZMK8BcJwFAfodQNV8WVeE4BZcemLpy6yoyUDDEZEW7tVhJZS8oHWOwKYe
yiHxBWseuJ1pyq6Pe/ucHzXP5JziagxdbiRI9sAiIx7h1CWfXPhPZcRKROjQ
ufPLYejzZbTkK2Z66TBk7TOJTQM+4ZlTcbXJEZMlrW2bMEOixq0dN3fVpql4
jHAoz8bAQBX/MSo+4dxV8AacghQukWDKiaf4Nk5h9grAV3rx27qHerxwwChd
EPjFbQgbJnPBiM+yxPcqjBIN3xFhqwN6A4Y7tpC4H1QNCIgrgknqWujXNduW
foU2W5wlCrHLKBRYXYG9AQqT4C9cT60yXxmzslot2aBNT1ZiBiSxHKnQ2gYW
wNz4r6bFkCMwE+JobBXRmPkludwrt9mIakcJIRe2oh0SPovdmhgn2d3Q/+st
KiVw1yvPIP5Kito3MYapAomaCX2NCwtL43oIC+HdJYY6vh06BeJKZ3oE4uxZ
TY4RL4Ubyf4HIvCBQKioUL9lz+v7XLaZDqYG531voDJb/3do2yyih6qy5Cc6
NFTHGNe10yMvjRg9/zPa6TzFFWQVP+4Bdk8RD85ttFHJhw3Q6Rm0f8H87C7d
Mi/a1mo5G566x/VhK4o878qwgmVWa1dihlJ8Pz0bdIE+6NKBzjGWe78LKqTq
KD/AF6HSnwzyCu7n/Nkj/yPGtb+6t/ScBknPzW/07yEQpzRki7FZvome9ZnD
gaipy0b6CN7KEwqsRSd0p5+XYBvpBGcDJZdsngHUiKyLTKhTdkkMJXw7iXhe
CNyfREe3O3IWGeq0wy8O1azpdNcZi8GQoy3rQcKY946JfRutfCpLAsozc5Dr
pmLe6MorSjjI8e+/ezibRXUPGMRUPNaTxs1/lEbJsncyMBA87hlzRAB8dMrT
ocSuemFYcTDn9clydUoijm331sY8shtNP/YG/oehF6QtjlaZqCcXuLLHldjU
S1gvAcvozefrWeOFiS3AtwxluPKlDo4hW8oYkN2fhSc11FNrJLl6yG/m/G46
c6Udk9AbtzjmW9HkWnnz4pNBsiudnCbrsgBZMdMP1L1gavbGzwv0Ol+YhvLq
B+9yc/ox6yIVRf9aO9Hjn8uOJv4NHHswUACAUJ/KfhbZw/HFzqdRvvshenAc
oMkXVkaeIjiLrCjogd0UT1ZHU/4kFqpXuz6dlUeMr34jwq1imFWKTIGQlQSp
lo8YeedUvRi3Z+3nE1yqwgms7BdVXCuGrlvoitsgCkhdxHlHNZGmeheC9Gmn
cg5JQd8NpntEAhh8AIsafjrKvkNjSgRyaVrhzKtuPe472YwXiGIIUPCbbx+a
UP2qb3Hf22RTl6RaqWFurCrgJ75H4kfR0oJfdRp8QDKwJ4sGe+ZTnPMrBi/f
ReevrEOPgjYrE2TrV/b9YeJVu2Xsjq51Gnqjw9m+LvwsQ67GYv/4GcTJ6stn
ju6BJZailrSGpdsDMPkDzW6oy4ssaTYHSvLHTL39jUp2ykXbbCftp5V658B8
Bj+DytV3V8yWqfrMZAWrwAu8xCEPiceqEDZrTgR2OoyizUNchyZl/9J2FitD
RPfzMSI8kJhGvrDMmOslwoSBv7ayf4xGauWuHYw91T5HUirMW5RYIRWffV52
rL3hG1PYI8CSxN3JRKvBNqSJsR0OFL7ETM2LeLgpOGqfkN8LqY/gKpj+uQoY
LKB9Rqv1YqiMqgxB9HPKNVKbA/ZEilDIK2kga/2M+uaf5ror0fSGqsOsTaZb
jYLwLUIINgSW6HkjIk7WNy3in4EEB2pbvPeRZSMO29AUl5x9b/GUaE0Nh8tx
GYv8LrETkOSIIa80mHsRNgnRoFDoqgNqAFe5zz4WFrqci+ID4wqThRIj+KSs
kzUkkdtOtq3diMrWsNCkjve9Rs9I0cDZGt0zlVZdVnJILNn+y5YnlvjL0TYY
n+IHCuF2g7ydlehiiAD2x8AbmnTkvkDGvV2sCT3pclWQ3bI7CuOnHCeKXYLv
Mo70CEBwcY7D4lc96CC6L1vEcA+kccdfzOBZN2XZXK3pjQbOZNUSa3o2wg62
J+kEkOjtF6oeLDn8ipHO0wJZShbdAqcIgktig6EJz7vihTRY+ZelOT93DVpg
MqsN+fUQFT9oNxEcGJIvMJj9yp6KfPA++AfHFbkTezd98rYX4mMwD1kzUvQ1
Fa2m2UtgseWKBc6AIdvDMAH6yBCZm83/vYhcww0H47O1pN90bYaBW/dXQ0Mn
mChaK5j2RMubpzh7f2QmVcfDVdZc+yvlzslLOkNuRKsB1Z1WjOqRM4IBYDOI
6gM4TPspXKaYvHP9w3ec7x1QHyKyvfqHfm52zNiiwfxDBmMFc8xgl9wOUWRU
Iy80E8CCI7C0pS+ddePxInY/RpYeZ7fP61QEbXtagZgrZYQsi5YbQV1kbTqG
6cBoQ6m8+tFGnyp/5DArWUxHJRG8my0zDd2uHdBGj3b4XSn85hs9euZ0N7zx
ksJZWPe0iseSNKdEOy+Z1KsT6ms1K4L5WmitWvBbvHB/axBTooTI4vCsvQXI
oQ251C16TH62v31EVD8ABnGxILgsuQqQJKuEmOfeeJ5l5a7yQoJDRLe+9qYA
jU5z+KpGlO0OPe/cJ1OXnarkUjHHUb4MWMqm2hLyucsI8iKqLS0Un5WPS13B
oQX1Osvm+pIpO7fKx3uNxP7uOlNuTCwWAgW0pFCwTcalJfBadXHytAwBnwSX
gfluXZ/pFuY+gwZ5TzCXMFSBBdzrRNS0ZdjYect6K/KqDqLsye5oHQ6z1Q2A
6LUY8HgVVF3cRj2VASxkh/Ese1FvMeqRzej+CJxl7kUEVvyx3mUTIY64dXht
iKPt0En/70M0v6cqESqAgaR2xoua/GxmqeZV194FDuUiLlFd6PCHgHXOJwga
Mh9sq84rATPDz0tM8v0TXyjOIwqlQn1MexZ/9kmMr00IePtFjObVqwtfUEEF
uZM36kmuwWQ7qBkLv8frY7kHqZsgMNLYTaRbgA9B9vm/yFer5bVlt7uUeLmO
HirXlxgzDlE2cI+MoJrK/GDPBHadnkFTFmKEWHmyxplHhIT1VgPuLpQIKSNp
nZDtbgUWUVPG1X+7HViqQcwLzzU/uQY+9TTz3SYgIjpmOPBc+q/TEh8ROg6X
TKdweAKLc7N4oE4v3cjYj9AsTA3IRhWKU46hGgLzZ4kbWIAMADtYAlaWddFf
PbW3v1JU02kM7PUwao7XwXWR/Mc+0KD/ScspBxY12oKa1mslD2NPT/L5fpTK
nLpcfHqlWygFsMqHMhl5egV4P32oBreAM3b/jdjen5+YCfMv5U8z7XPTfnNE
oUSo0X6U24zJmdEyNLTV3T8SZsOWHa7AUPEtOLjqD3qKqg1DvSA1n5Iwgwye
L8gGv5Znox/Q5oF6QC+sudgagi5buH3YWZqxFa9c9k9Tne5ZDEc0zdRgtheS
f8DZRGhKds81TLHtbU1cXR5atuEIlk6aGwjb6IZASuXEjbP3P49ijKeVhP+S
ehLiD8r4zLtlhV4aJnFPxxDibGCdMJ/dEPY/s297dImYq0YHtV/cXE7IBxm1
m19m+j7qdH+7oV+9gPGOSmo4/yV/zC5pJf3Rlf0n9DXDlFp+Ms8NHpTQPBMo
QriKQAk2s7ZwPZMiMWoVFYEk8YJHUg05BZhBeV/qUevJl300QBJBK3fjKSpE
cvLzBQK7P8oAcYamDlHJAMXQO6NKZOb+IbLQ+uj1kdEt/87SLlIjrGE23bDb
+X1HEy0l8M4r1o+FgmB0jkNDPBp0U3BoTJgS/YJL1TZxqBmFrKMczETO3Emg
Uw6QzRfYLbOYVOribKAKgxHkjDsCHzrzZnaZ+0jX+m7y9N1o8q0+hx9fz5fC
I9BBCWrHvq9rjaj9zueavY1aKPBaPIzyURHssg+xg+DwnS6/UEaiAjldo20q
E+I5unUWgw9SH4qxgGSJCl10aAVD/SRQL2mux6avknQwbrSSlmQUuW95i34y
2JCUTTX2/cyTuwT0tEVbXSi7PPj0dzCiq3xofj48gC0hcriWv51wySDQtd7t
TCogBjJCPojvRHgM9k9m2iGwUkPq1NoH6ow/rFfv/lzkjkWYEvkoCksUucEk
W/tn4wrRhHMhbY+1Kiil23MmZA8mVATDdmQw+kB745i13Yh88+AMD0sxNVt4
4d4as2hfoK9evmZ/WZ41ubdOxKwOPLP3X5qxcH7tXVRd/2lRu6CqBy7MgZDE
MZTo85g6gBB6mVwJ/p3L48WlhgkGKOjR54BM86u6S9+lUAtJG549n3Ze9wIP
HduNfODOK+VBBTHr1gh5RmxrUYroL/UsrXRImqHbhiIJArL0F3aobXZS4Hmw
1cBwr8NT/rTRlSaXvvFhmHHksftW55SB+pdHGnut35xg+absj3GKOBVE3ePb
/fKpzM1HarF5qk1IH3dfC1OzHWC0Ve6NnihG+rT550bdqQMOZABSnIHr0/xU
d0ixSC79B0sv5QIvA/tMpn1Xqk+0XCWQBvUvMsaKdd/0WwJ1r3YtrH3iWWPQ
nXlM1x8GHW/TziOQGccpNlnwjn9ZtUaB7PvBcqFLdu/fgpucAwAaP4N/b11K
fXSdEwBrnxoU/5gKTQLisFwDaDmMG3wpP+GQeyDmiTsEuEteQdmvEUlg8tHW
BvJpveTIayyIeRc/QrQRMxj6zfnsWzmGRChCNHl+rjtWhS1Dg3P2cXzfNaV5
JVaix9CinjUTGUPH/2nAuc76T27Hm1onrll//6pan53zaU/EpxBw8DixJoJv
pOG1p0vOVMC5jk6BOiRL3oJqIHaejvkd/YgOsYvE5L307hAIqU/o4nCoVR7j
f2PO1TiAcGa0fkWHmXrwSzRMjo8+V0hEs9HQb9TvxYqEjOooLwudIarjS0fS
+WbQ88xI5kiaK+MVxat3JQz3LGOm7pOaHDfvAP2R7B6LBBSD1+erpIo5wLLt
NaluWucPrE5+6mrMRelHMZoolsHdP+5DmlQMbGUMWuUKs2dERgd3Ev/twz69
ZNhXqqWcc0ihbtZWLBa5MjGNqPcBGXaB6tlnxuADRP4dBLmCu3BY3h1YW3sh
ZOqw/oENW09kuWFSqGo0dn4iEdyUwIN0odTKJKqi/cKVYPEga1fmFRiMPirm
6KkY8CKf8LNFfxMIxSQFKOfwMbs7D7ZYR02OtoHOPFG5faiSS3j9QiKmvfmV
R74mJ0hcfW+okM/aW/nqE9RJx85UKQI6X/AZnUfTZjFyPBjm/2f4roeqjcpY
7UxHSkLuivBxluYexJPzRXhYJForOi3bRooomJcO79Viac1LHz3L+SnSyWm6
j/Rw/faHO4GlfFKZZluHtgs/kLDAdzC5JV672aXp5BkbDwDHBjy5C6swkfNU
9V85jG1fZ5nxD7gyPjUEMhIAKhWjc+Ii1JdHgz+XdCwCrLZdCH6VL4axFvdj
1B4ydX20m0Rn9xSK1LyUS4FT4eVx0E0OUlrJnCg76NQ+pcYB65uuHYITkMKi
IvVqr3ZoCZ3lQ3yi7OwPZs3zabAcDO+0KnIOANWq/9pkRNStBEj5iT9YHbBW
igPrYVbZNtjhHkLVyQyPlqAP1oCMndzeXcYckqZtxf56R1j8scBoHaTvj7tD
bJ951YZTJRDL6mslrKmjg6hOxWXg18jOt1bGVI1VIuVxk1SWzhIn6hvbIDvd
1GHyqDGnOFszAsqIVyMRWXq80OjJshdciMZ4UgKACcj+xqQzaNQ67C6QTEtv
2eQBPyUQpJe7QJ6QUO8KgbUPR+w8RGnyaQDFLyNOlxuqe3dvW36NBN/Nd/w4
iG0NZkkHTGvLKg6yccgrNoUr5ZTaF/NwoQkwrrSKV46lMD0nKlVPJNhq3W2K
MlWCCXvzOllMSvJFJZdszJDGdI8AGiB7FFECunYHLEOTAtyXu01nAkHaKgpA
oaI0cpnWn3F00cH0LdkcqtxR/sqbweqyT1hcyicz98sNRHO1Ea6DjFzQ3ecw
Ove6j9mHpSf8I2V1n4c4WkxTbKV2GLq4Ov6mHPeW1yt55yJL+yay5RdbpZ4t
7KLPPTHrqK21gWD5JGm30qydBPifL30XNe7qdi7qMa90HXJhtlx5rqBfqyfl
mIkdH9VsyonxNKulOxa9xLMJI2+7S7qlO2vayH4RVbsTF22DtKDi9pylqdio
nv/Eka1g8Z+/WBYC60vaWmaF9SfvWXflRTDSvpEBlY9h+h30ZhmW+O9mt9gR
Zlfpvm6HoS0w753He5UrfUlOkDn0OJBf+Ca7H+5UiL/7dd6AeqKVN2E4/P6A
5IKu8qpTqKu5wQkelEba9cgEYbFOUf2hyJphCUj5J1vpIkiFeQ7iaMc9BK8a
dCCHW3xZyXr3N/54pdmJcoqMJjeEn8bP/cgH52ipDHShwNfRqT1JMeE7HvVJ
81SXh5j8JuHRgV53dyGZMd8uL0kyIEEu/kGaMyunsdscNnM+z1HrcHceOof5
0atm/7OWYJZ3zb9E0wTqiSs7MRzB3SCu/qwCrt56mxFJS8Yj0QBeDZwjVxhU
4YWEK0qmviZB2z3hUYPaMvkpCXNlw70TJh2vgVh7cbHQiThUw8XdruqFBl3P
pzPrsgUQ4Z4Har5VTgf1O039cwKOZN43nPjw1lop7ECoZgBNuuOFjQBAgjgq
u7+oOTuf1i+8ZqgCT556hOZjuSv8p/HOu7dVu+WhXk22mrRpDy7mffjcNdMO
fppm0dPLM5VMruQdz/x3T/ab0Vqa5bWDPYgfJRNOFx3duu75KK0adNkHYIXP
Tm095cTYnqa+IqTZNHqW/cPRIofJAer00uz5NHyossvSX8hTbuWeRCIjGkJf
HCxojnzFuElq62OaQjfUX8PJEZr50+JZlr0cfJdWcxZRsszLiP/a++6l7uvq
XSsx6dj6pN8YAFFRnDz0x7aiYT9R0ZY2FHbkWvj9/mp0g8HtbPK5DFcsfxEl
00IYwmtCarpH8TC9mO+dqdXEpXymW9m3GxAW78KIoBy+Y3DaFieIXvRVOqs+
B1AFbyu1UEgFXHcZSF7opD8ULviYBJkfDaec2K1gGX94h2lhR3iBUVgyqRPe
TXq1x5jWkmGjDHyuTA9Uaw4OA2oA+kafKgVJyo4T+bmc6HC/JeG8jW2HHwqy
JfHxl6eqGU8ZHGv+MjNzAUJyyTVMSLdUa7Lh3OP6nq9n8Qz/fqDs0YShnQUE
ZJ4qT+IMwy264jzfdG85/1N50m1APHD3FZ0ZXO4EUn4m4JYOCNAnSLxtsj5U
eNxTH8gT7Y2s3lXS1595dG3f5Qv1jZ05urT1sPm5X3GGBcwqrAcdVCzQq3eR
pQMO3s9ahvtVRemqh4ACVOFeBrN9woHmSDXJKpxSTUja7PXSGSSYTgalYc8Y
9eP8EJtvhmlgQpEA5/73xYmaMFwX4UFE1K0wyzpoL7+W2A4vnVnpHsbG3Mft
ZBQnmbA8Sqo79EUhIx1AYS0/cu5YIjGMmZ91xWPiyuPVjJVxwgKxY+VqDnRb
YPKVgEi68De7qB11X0yRLmzVdlpySZRWJBDV191FhRtGGpp/ZB3CaMaRJC2a
X40XHv+VLluKEZim/+O6UGgqfmR2DuOHcf4iEPXSDNEP3skMMf7m3mX833fO
CvWj6zALMhCr57kxDIiLbAVH0tVbXcEYKTAWeGrZgCLnUaQQSdC2/TMjexN4
v+oBw4qD0c++zqm6P74pPypRsuB+eAkv22wOcaGRLv8IiKSbs1095YsesA0M
Ze3BXEb/VROgDMjiij5MUzUJ59cgAx753OXQPEz4tQIzAyZn+oj5xUGNo3KT
BVcDKdepYeNDjYE8O3WRoZC6Iuj5NE+WAExf1MsiQQJSTcrmjcTDIhJS5wCi
8UA29D7WPPLWlTnIuw8XiyNwawuGC3zg8g2xp7vAu5GmdVC+DXGg6t7CnIOa
TOUvc/Pj+U5POgsPIjnESphqSPcDuBOQTTHrdrCLuuPNPI073ldi3LtBWHLu
SywPYu363mgFkL0q6xKvnehYhlnH4UZ/gQWLCycmk3GX6WUKq05gwzqerici
utVMUyvpgBeoV/8nIst/mkY91j6rKzHisz9+9ukxPdHtn4PryKZOsaYhJRhx
v6staSzQ4z7z+v48vPaSc5Qho/2NuElI38Zof/TkAfX+LymsQYBrzmjFHhYF
Rj1OaoCUQsex+H2EqioUM0R7BdjWZc9jnOpes3Es8ktrCpfsvNZ8nXYadUcL
H9Jrvx4OUwo7kI3huu9ITiFVwEfo7cApECMjdp4WPpPJQMZdVteeZgsHMawQ
OrT0JdhosTpTDWEF8RJqbB99ou0pnbkjPkBud9iNCAGFFz3PuyLAv/yVEbPs
6JaYayYu5TlNlkdMmmm3DMw3PRd27W7V4EuKc1n3GckeAkR/lzIM9lcSrzou
9LAX/1oGYo9JMihM55d2YkXt7sRUef0xBdjo7p82ZnmW7jJvTAvV1ySJdsH+
YhEAGL1V4T5IJ98irffDYSV+p7Upi727g04laXAv30Q8XLDxIcmiWgKO1ASP
GsSJ9+PiR5GAx+IhVeAPS5NzdXv3E1Sy3GCxjbrwtNP3j+cLXXck0LRRCCZ2
QqHymfAgdHGmmtFjwdbFnUJOxpd0XDULbspShZ3t9SFQdz/aL/zfJ/TZ4IQi
vi9hkUfxBxCNSL/UFOdnkufFq+6UXH1QTU/ppq2bb1Qlc8lic03o9fqQ1oJu
9kqWMaWAPgfzYDoFmzzUH6YpWGY3T9W8P8TFSGe2oU6wYH8Ib39xQqwNAt+a
SlI4fbrBFD3AywSCLLAhbLuUkhngItkmKNPbEQ6INnLunMKzhMt9c0lKirow
vMcLjVRPb0WBMS2++kbkVxS+eo6eKHjZz9yr97MOsotplS1TZX+AglBOZlqp
0O6hDVg6yUmVJ9Fk0NxxDyiPbipR82E//t+oopjSfNUQvCwttWHi4G6X//zD
GlXzrpCO6vyalkCyQoI/vhNW+2fQc05Juj5Rc9X73ssAGyw/NdcEdDQjC+Hi
ibqFMpkEckW69j4KIjTE27tPi4mvAD3NrVu3+PpdGxP9BqT6Bvr/+odgOcyF
1Iv8qz8cRncsmWnZOxmuGKDEYd+Xks4+pWS30/TxS1Hqoq1hg160kRj4ngt+
A59HzLxTCIEfB9yOy+wlYVMJ8K6sbLUG3xDX1VbZM7OZtOoLZbMjaOIXaGPC
hU8itt1URLOMi9anSD1D0b5qPay6bFe0qkb7o2T3U+P4y3tY9w82wZbwLUyy
hrrBcr24upwP9oXIUWurtQCGIb1ZFG5IX3YWHusthR6UYvL8zasyVrdcyOm4
5rJeUwtlQ4Uu0XRSkp4MBm6x8odgfQJSvyF2D1s+kcGg3a1e7LtPJ8eueFFF
vwkrlIlzbFLy2g4spRebXzCnDDVZGds0qXs7RLvLTqnoyOneP6RZ3FznDnoK
eEgl/o/6h0DuhVcir/DKT8CciiwxDph8sLARDn8mZc51o/U6Qu2MgQG/sn4Z
3RzihNUml8zj+BsXzHxjxpmZ1FSAbmKmd+DK4nH8vQIkKVDmkDM9FC2JwTYM
dJXkllj/YrVQXQujP9mqCN61ASLUqjJg1KsZgdbjL6kpNZ+JHVvUCX300OER
/U/HwEmodB+kokFHVdokdIjubgTBUNICnhtA/CYfk1OMPMQOg5CldJh1oHtV
8WOqdOZtm9iaDhKXZO7zAk/WyYMYM6jfBwy3J2RuZTS2+ssJIFjs2QIvNBSM
eQSF+WfaEhVgyJZnTphWXlhrzfmoNRUnsGW9wsxRIsjZzlGwU80IUwaCDLCH
ZItzhYT5V4t/GQND+/GaxR4d4ACJ/v6drpq5zY9iGP3IbouDO8putUH78lKr
tV2KVsVr1XUQDB8Cu6gamyrgri67H5GUhoethd0voJsHbS7abXPJLOzHgfG/
NkmfvHrKTvTRc5rFbQcvlG3D/OSHmOqQsQZE7MhKpXgCS3ymplnoGLsswuBc
CX0B4z+r1x7IYSu6+Taa3bdg4XIZ2gTnyUDsH1flwwQYmI5zsiNfaPZjtxSU
UWlbDSiqraXCRJR0eTomhbJD7SnjXB5AxeMWDRDjwWcTSbPr9xjRaSKxWkKf
dh6O3zi/EWQm2iOpkxlegyiqJa+mjTXVa/TC0CacbUClatFSlwhIq1sUDixZ
LIByFQ9T+gki+Q64GIihlFgClb8vW5Qa1qMBW5vH2o/tjHdfxSO6bGYd8OJg
lluTjIG1nRlO0axey0NS9eqSnXx0LzLEJUboDyXy+aQZra7giizJAc6Odc0z
jQvTYHcoVuL8MSxWZ3rTu0W22LlntIxFov0GVNSjMGsKO6lVc7CPEUODuA//
G9FnOHsnNfwIeSO35SPZ87pEtezeHu0ssq7d3Ct+jRucr0qyrAmebi3JFGON
Sd2esjRD+9/6l1ImnNyowNEONgTnbyE389+L2wcqUJyF71foz73LJexuyfTQ
/s0dcE7drXcdYXAHaaqDyPnUng3s2PEimGyZsWHxyroQPKr/PEYlPoFgB4fv
BnLSvYb4TmprjCicjgEdoL4LlttUweAbGN6O1Y055pFl5KRaDFoug783ERyh
U55Rb18xc5suCqHd4d/+082SsIouXDi7aAjt68HQqDz03xcvJcnvtpJ1Ey2K
O8on/4aKbs2jSeMBFX0dBY3jaPDsFYC3IGsMIBi/laAi6T/ZFGjAVqUFyRNZ
sDmU9g3Hu21kBsCV72zsvHsf3+8KSNkJJppj39lMxshN2jj9R0S2YCFncXsY
JaKtFYTYrUOwjvCWobPJH1mFi1luj5iAivnfJLvuzCPbS9r6efqBZK24HAHA
cYRrzm4mXz5N/cEYEW85hv1NfZp3Xf0k5wdWUQxkYFjLYND4/i2peM2hkeye
XvIZRnqbaBBzih/6SbN4r98/bXV0zGqgF/tFThWi8VxUkckNrbh1ktswKPC+
tAaHkshr2P6nOfUd9zJs6rDw0Pm2As5zSdHJLOr6T0AluRaPMAnhJoIh+GH5
AWmKe9+mk5a4xi6UaY1PsoJ2jO4hanOwG3XWRkQamsswQyw5eW1Ejz83f6fg
0HmBxB2Jgip5xbhJSuJ1Tbu0c2ZoMHRxFZkzfF0Qivw5EPZua4srZpLTFpfT
qDdI5eGV9cuiCHW3fRnsTC+uQVF3ETH7zB60HaSGfqOZe0QMYykNAaDiYmfC
K5UaL/j+adUdqB2UyOZTQXz2DKx95zdia63zW0qWpJEFXM+L+XreE63FbGO9
okOw16kKYyZIsReNQD9LnGJF+xnz7vHp594EIN5nXB6HNMjtJiLc8UN6Wf1F
+BJ/Q78tYGZtWo+eNSSSGEiM2d2yWz6SVDK4+QN8mNPjBnh9aBHPpkP6aMn2
CVx+h9TERiqTC/D2WaGsqHqR+6bOfHfCsuqVqOyg9IPjM1gnXGY6z7CVmUDH
cVn9EkXmELbDZr5bfFyclZCSifsZmxE3DO5Xj0l/gbQPgAqhTflNUktEU7QC
EV5+vTHDb/JK3iEihdXLOHYGdAZauaDX/4u62moVcpB7BMwdUeGWZM14mbHe
rGpFxVxyTE0CSbs6zyfZL1Ju4Gmece6JwhvWSUGKvqGYXpaXlDh+cx6vgDJe
gs9nGyPnl5ByJkyUzcu95nTzHa2JydbtBd3jMZxdN5bFA/EVRZuMFdMi1HRI
yOjgRZTjwn03WzZ6tVzy26JndJ1IwEyD6xZKCJ+i6NGTX63HshzJ0FIwwTAd
Hp6YHh6cn+/dA/G8uokEbAZLLD14OUXEPdGp2Ep3yJpX04Nc6PatHNT7vX5N
phqWnZ5p5uH5iy+uEPlaN95kcq84jxkaydmqhWqTfxGrcDCYIpW3MzFgL5cU
REWT7goqWxuDgamhmZbbHeu8z+CdELejQmAvGhEghxfY399en9UbP90hWGge
mIeIimN7iItAlAv3qLbNDFavm9uGrQRkykSLvMKyX/PdCf0o32ETjXrxpEkc
SPkZRskQSEEgnqzY/OfhsMLI5Hmx4hkHymueSNqNf/4fDMyW9Utm0JJE1S3o
fNs+2YE2Zw+iE/FB3ip6pX27mmw/9UGBmnMZD6v9XfEyhENVwKXYD8nmeiIT
9etwUpC8kflWrw4ZBMinn/ArcYwUUxHWCoKynQBtJeE/NuGcnMDC5qfkuhUq
ID+L9EQGikmbbOyAjVK9/uS4nZKJPXFbpTABVtydcb2bMyYOSHOCmv8Jqok+
+3fZf3StrOcUO46D3sj2ZiLppUwJVKSPn+x4E4dRVZ10fXcojDf19omWfNOF
taL2Um8d80oCQirH1KT5hRdlF/fYFcjFMSfCuz2HskdiuBOyjIjlTI7Qs9PQ
h5TdHf73iKSJf8CYkNDMx1yOXv3uLPC69I2LuyS/VGbnaUFWNr+e903rHHSF
YMMaVpplI7QCa3qFJJwKiGCSxDqWWk2JHXU2be2vfjLTK5c927eRxeEEit0q
ywLU2pAfN5fgGHjAFPE29RLTKvw8a0B6WzDpHmBI/U9nSdXtu/3CkHoUf6YL
AuxDetdnYL6PGELZNhvvekpykz3w4cU5dSY8Fc4TJUpD/Rv0ueKzR20zVhqw
AI7OFaKRe0ByOSDEQFRoEWUmCMcjCOk4ky6GE2kjITYiMCOGIUAkloOmtZAQ
O6XkGG+T+VcZ+P9im8kVSmBrj/rvoegbXFWRHTNokVkJxGAcvcpPkug8htGX
tMSXNjsBdBAoIFRPhDIv9sWXwhuclczqqCejJXVBk/duUbAAaD2Ci5G41Cmi
/jFeRLQYluXUJm/l1K/REcrVpFlknyDnVkEQzr57Qpck3UdeodGAMZQyk5SW
lD/9cMrdwEjWz3zpkFBlPllIRrJj/K0orVZw+MvGfn4iEukve9BJ5cvugyX0
BhRX+NcBHSFtoSJSi62HrNuKhwRVqwm0Nai+uSnkZt5BlXALklsRXRLBkO1v
AgWebHAj/9dJdXIOuTngkMaE5UEapyRkUwxnw8bhdogKHedhEuo3F/rZMnvd
eUaykJ1Ndbmx4Eg9WPL91SncWepqEePAXQDcUQ+dH/eq3wKoyKwtgZCC5b38
rtWwJheTxTQv5SnO+JDWVGQIsPh/m8FozebQQ+n33vxsEKNqsxKfJyQznp1i
nnAgAqa9tZECloUvkFHzn49Z0e+y2NoLz9AILkT5yWn29i03Es0lZzcZm8Yx
Fbe0ZkAGzjEil4JWWUNtKSPlQ5MsynD+weva5uD1AIPHfGZ7lWuTmyuu0dyI
z7kCKGoeP/+FT6uOp4IXM8WuTYJncdpxSnpR0uY/n3ddhEiF7VVAhmWwghGz
0XwQ+fP+qtsKOsERYVkIC6YRbq3+ar1HzDEqmN6MP4neKo0a2mDeYEiUxMPq
kyGL3nl6akKw5eZ3kyZKZZ4fpVtDMb5kEy+Avq9KeUNJAEb9a56lIjm0HLnP
f+HC7yqlwB4Gcmp2Y6yajDHpzfxSBvq1/mknHje+bRznW6Si4UJuDi4K5hQc
e1bRRyQG2ZeTb6g/i0Nl9BMXbuK+fSy5uyfWAfDeyInPTyiJXkQ9F+0vNOAH
2dyGCJW5p0rdLnSdw0ZWyzhyHxtpY2295jEX21Vvp0gsB5q7nuXH+Rs/HjAT
S54cQ+axG75nxmN9+EikaJxko0w8s6kJZNs1rx/i6D7LsHaTxlM8kz3LmdQv
xuYCuapLWcxs1AwYE1xhki7uXcmmiX7dA2T0bAYYcQfSLeutNqLi3Ceh+spA
V00iA8+2UlVjtr0D9bxJPTfq+k0wa44Ib/GZEpuAMH4Yt91WSuIgU32Wl4Om
zVah69DKOQOVL1xM00AVPDGlLi42C5YOEARdLiRw1zt2/v9p3WGqz/yqY3p8
s5B01zw6t3/pUb8sdNmag1yTYDXg/DNekYp9OGEQGh7aiCmiBnS44KyW5PhH
StRS+7QL481csNdj55yE+4+8H1OZHd2ZYchZdKKWCr8JOvhz0Rp/OVosjnWn
DUOT2c0khmk9ojNhF8su0HCkxDN4Dj5lwpwycPMqs4jtrFaLZxoCYuT+qQ5I
JasAiit7gbODwvwwMTczdM9FmBV0xdMmUxs4WqOk7nOLGXTWwleqphdVgWh8
VWGT3omu/3SMCeZvjF7mtEaIrQ4g6dR4gVApyhmJI4gmdsOUmWDWsoCZALyY
/lj3qe87H84u4GJylX8kdlEJsk3aoo/Yhp7qDXfu+SF+pCChpPeUHIevSE7k
3t0BX/VYx1qDhUjVeNkhUBn2ijXwIbZsfmn7F8dCCX42MSemyXnZJEixmGOm
LPHGYjMPcIgb5ZjLvZFgFdgUIKJujfdtg9hmeWVzrhp7h46mXahcAU1E/1/L
E8Mtd+XjBWPEyKD0L736o+oPnqMwcxd1/6sSNIGcz4L8dy1HoJ0um1lu5inU
Nr5MECjeTi+x3PxB7ltdjLlqxFnb9mraQ4Ev5r0EVPhuFu5yGe7R8MhqQ4Ln
WyEmBQaVP7A0oSOokBAVCO6Mge0+DmR/TzqjXjQye1Re0A2HNfXOEA/FG7Gv
PrggGKSO/6UHN0SD7E7YBgxB5omgIEoeb1fVlxbP6iNQlUR+CgeIp3TbttHz
XPilJk0cVGc6ScHAgSuy/gtKAp+pPrWeiCMV0c6V2lkXIgJ8k1m/dFWGBwPh
8bZHm8OVmEi7EqGbmRJ20pZgj8CF5ndDK2yPJSuJP79kz4gNmbsmSmxBm/FX
P9q9HsnNYvvgi9IlTgU5ELEk2ouOHnFC/G9akEXU+ajg06vwgKdce/oYS5LX
2LKDNlcTXCONli4e1UcaFlrsePJgzt+TA32bCqiPYMeNjcXU554QS4f2BPp7
5jQ5yd3mJ1+LR01EujFtOWnCbym11nVHPRzlJdZpGU/PenwYm9+InBtK+iTx
zzbEcqDQlVRTG0k7f11raDzUGR7lbqnX0kw3XQcdau+rzUociQ6pQzMg+xT8
WWhPOBT6x+e8N4YSeEVwZW5j3pCTPbYeXh3yJcKg/pFcMgYtXlUX2TRvAhMu
NecZJP6v25aylE7twDV7vPpGMwZ9a+JudYMWC3/uwAmqtPD1joyYxidoVBp4
XUTAjnvOWab5kOIDrsuIHkdgQTP6nnlDk35ZZ6RFSzObZ8YpPe+kEtoQkyZa
RLBv/JNHOe7SFOIDS+TwxYOYyK3zUVQiRaURZQdsZGT9d3wZ1kbrR+JplZIB
qWAjSEvxhoKb//3YljccVpgP3jHGAFhO5XBrzNt/4kCajsSwALg60vXc8r2b
zG5ZGeQ4+Q+ZCmzft78YG5xw5e/ZTv6zZg4TtvXChU4fxYA+CIjPA2JX3QDF
dzpgcTj8GkYi0Pl8kfIMuLRIKZjvGPZ+8w+QM3gWb6xuPSRJTK3mqur4qBx5
gb5pPL9h7J5AVUjcI6KiWDqDH0D8jPtxV3nyofSjA7/lqGRJ7yQrMIAqs1Y7
BhfK3pxDmDeP2iANowo+W4Oi3CK/05BX/DZRHMC070rtx5miDlCRZxY6Of8r
oj9Aci4Dd9J1lOU+QoJ4maCXP40pPF0gzGnZ8KBkGAeGsmgmXydyiLLBtrxv
St2Awn2scelQo6KsuR8nVrQaifMNDr7Znj8hzyevE3DzHqSQRFyL5O77FZH0
n3LDI157lYyCgGSLd+P6u1riYPnDCEZ2CsEcayI/qgBQWWSTFkIx5oiik1BY
pZtE2PcFzVq+6Su6QO7+hUVnyPtO/OQis2TU0l/idd12Z2FUPWRipQCh3riR
SD4BDPkQIHZbhUdI9qxpmmRV6NWnu/XANxWk0TdCjy/u7Lst6uoS9ckZqxJc
RzBDlBNqg1teH+lequPe3O/p7bLEqj3x3w9kTNIWqsWgL4avFVSHy8GE7x87
3G3V99QiaujNkzlhlKrpeqO8SYczsCkJFhNg5mbcBzMfauapZ1l9SXPNqhmq
UjfwW7CrPTbPU5tO6S4V5N8HCnxlUxddkpkfeZ6r6sXAuXfwhQyO6D5H52P0
pIsUd3tNlwvYKXDfCzhxSa58eXepdKYM6NtzvD7jpARbQ12xHIs7A5kHwk7Z
U69zQAJ4j5ZASDOk5gqAZE9nCynmy1+BA36bt9d5KwvgSvn/yFVvh5Ekj8nU
8NrPC0R/ZRZSP4ibE6RoFhYQ/GSo8UtVH9byDBZazjYkG3rdx3Q78q6/3WhE
9HVuvcTHd8TeXhOfYVnRO7guCno7eIbc5Agpc/NgLKsTJuoOwrvN14Ydur6k
puQLb9TNxyj6V8xudmiz0F6ATXBHJjp20GTcD1/OsndZdTThXk4U80dl8XWb
TO+Ahdt4DutO5bor46/0zLBRjghmmQQhPYuGlp9lcWtZho4E0Is74o3xe50q
g2P05ly4wBJP0SIAl0ofFnxWc73okUS0ijeFqP5OIttAqcu4SV1t911HItfE
KXAJQdrArwhbrAs/majbmkQTHDWJ2VSY3As+m6mapELY2jZ7f4SORNXkaaBJ
AhEhXU/A8dfy8aqIQ9O6oYAyK3xif5ud99leaUv+4j2jjV3Wmfo9XG2U9Mnc
jmoxM12/xoqmCQAo5wztYnrGbNLPgP7vag6KHXwWetVj758rm+HwWGgQisyn
c0hJM+PoRm3HPHaTSlhIeoX3lt36QcgqrQJWWCEo/DSIIdM7o21LFcY8RulI
A7pOQrusdPkJnQ41tNH6s5n78R9JHP6joCABw6433QWUvI0yIl3xEfXT2A/n
rcZ4mNkeqeDATY+8abUvdabsMMQ8lzk7dUN1PeB9cXhW0Gq8bCoYOBQWaQ4B
Hkoyu1SOEK+BbsJdg1j8fCu8Q0jILF1RL7VSaDYIQDVpz1MG45slQW1Vsffj
1ihuB/fPknq0UYtiYbvio7Iir5Lih/2NhxooETHUmxkCAwrzVb1H8nyKgucF
U5sXOPRyKWtoII074a7X+okY4gHJEj0N+Pbnz1mtyxVsm2LkS7AkVnEsZT/R
wYLhyhrxgYWn7nRAtregAH1YdmuAfUlQZcaIt/j8vIuLAhtENdWTjwyXmJws
0b7L/CMoLRkJ7iskuahCSTJf+eHOh9GwEeV06vmZRjp7fXQjOADkfjYCpkEk
eVveDgWI1FKH0eOHvyjpKfhbTdqUEIjZq4ebCYLcHzu5NZL4z7rLDtNEftUZ
mexTip8fb6aWJoJGh7VvASQni/yGgqVoIxLmV/PZwh+gc2lPKw9EhQ8KXR0i
8iQaUkrccn0Ruzn9PKkC/gljV/DkAiuNzorxmhrzVc7O5TwtA+MUegEzBNCv
5Fa8dCVOla+b3HBH8VfDHcxDOD6XytAHVPmhbbSLHYa6f+Pua14aafqbg5bt
0r7asGRewwu21nrsw+InvVGUGyVMWyxhkvA5DipL649w5A7h1kWLjZkzIrR0
12JD1BdHhSO8IvIczq8WONLMDUEcc74MIShlXpqh03COxtAj4477k7oXusLe
ayznoObHUsF2LP60qKUiUTRkEVqBqgj8OJcsa6t+DPnLYkvgrZ3DE4UVd/3s
ncVP2SLPynO/wZs4eeDvrz/eBJhpsFl6KgWYInjX3RPmYQJCkV8+2ZqNKXO+
1548eU3y2f/E/QshkG8bhIcsJkT3JsrYLV0pnhyciVRjOBcX1fVb2B6a7Op6
3q+Ksf1vou5J0NiSEa8ylIne19cM77cmymQjYU7cav9Pb2JAE0PApM89znCJ
9c7yIam08pS8gG+vWES5feK6S0woTz+4049TxUgTresAEVXbgCarXxw9bxOK
oePJy63oi4BLZywaTDOxjhp0vum9kHRA3opSvvUdDBiljRc9ZVfABGfCWe4O
fdGmraJg2xQQP9EVafTHMe3KG+4O/2DGNEhP71EZV5wz8y8Sf6nhJtJl3mV1
g9D2IseqDMcPxewgC6SGaRtgQSEogdyFcCm5jJ9+pYy+CLdPI1MNYEVTxUq/
qEgVUt26Rk/B0hTjR2ws0XGrz8MOpgD4F5QDGq5LoRiaAgrnu3N66jVwS37w
NasNCdII/N65Clx/V9guTflrgUoswU8DeKe62KRKdOrCXVnZA2WiEv0L3xif
whOtETjwr7lSd/ij5EZ0WbD3/Yvd9RU3ICI5hd3W0qVx9GopRDxpFxSDvY+h
97nKnB9Dv/QoJYv4+8eTQC4Uq234v1eR59wgGDP7nBN1avCmpLCF8uCVmv+G
JDbRd6+OY1EYfN4amTB2t3c+7z9Ra6zttNYKHZBxI5ASbNUt3RHULuZ2eyzN
z2aA7DDboJ1kKtKdyhvuA3uAaHYLkSD5qOg/y7QKYjGxuSLnm7+iwUWbvaBT
axZ8IkmtRajJHTBKcyI9Bp/TfOeh7hwGowLRbjZOJdvcDdbS5fDKTAKtumIt
FoF2MDTC6+8ge7Ar+utEeTyXH+Zf3App+4K0HHkPOJi1/XYZ1YoRxry0OgzK
4jLzELxgrsT5/OAPeyffZc/yqO1RJ0JshBMXCk8gX15KpgTmUbQ0pp+1JHeA
Q7RX75tQoWK5UHYOHBRPK7EaJyiJjyGei5JKVzWcYyVWyWhnAqNhlhDVGrw1
ARUtjdfGofWyHi7lLWwA+bD177y/i3ASLRJOCt2xIsjcqJhnIUPpEUOCjAMn
x0AE1JD4wyMSYQhArwrbUl8I/rgec73TvdTje4J0bzv+qlVj3MsO4Vg4zJJB
M8CF0SS0psgSam1MqWgmo7/gvF8OgE+iX/GnQX+7ak1hDwZR8bddHq9VUd2+
l1lsKrHkRatPS4xB658+ZRrod02CFo97nhB+n/wQ35GTn49Lu1gQICIB5cs4
R/3mnKEgMxmQGegCmWGInjKtNlBjTpFHYNmV85gKopf2AY/w1oiEnxclH32n
+0dV4jkWelpHiilDRsZVyTWQTGxYrm/8WnJ1G0j6Tk2wAmGAbUMCBgD+UCP1
5pJmx3WbeDOI5t+1U/TL5yGLhU7lKVLHd0h9q5fAsIkkQbP4AIXB+HXofaTE
YSY8xQbkzu0ui6AYu+KiFQGaXIokIg6PxFzaR0rFRjtxcI+CRLeHGhAlu+A0
SoB2zUfJDfb6QPyFMBIZv2JSZUTHY52DHf5VPjIbjvm3e/MLkJSvVd+DJFqV
LQA+EX+yvGZNFoCJo7M+1Sqa9/nPe3U7c5hA7ssjUkQB6YyxF+aGbzwmIMuY
4LEdVQPNFMNfytnTOW87WT0BWEpV9q7JOmz+TtbmW9DsZooT6r/nl9LpSla7
fo2kncqy9AQ67XQ8g6KTfrvy/G/eUtF3pcg1xvT2nC0DvxggujvnQdEtImIh
VCblzDQ914j43cgOvwX+88pOG+MDAB2fvSrgiPvrs4JLUVPbo/VVsWBAUyyq
zZYkSkry+Nx1FX9gAdRrO16lUHGJi4nGlHsiM8R/4VD0zHzp3iI88bpF7TOv
C4Fw2HzixueHX27JnXKaKgcP6r9DCGVbuwur7N9L23IQaxDjdWuhabI2q+OY
zs9OSENH6BX/2ay65MgLqUV87ZM4NR+SpHJ3pQXV4Zq8q0dwzM4BSiqrF/nC
aNRLZnoDJe9B6Bo9Isf7bmRpePOndcPstqrAHsezh0LN1GOe7tbsGw73hEez
fSaUB0ezuFaflKWRqe9wZiLxbYnQPzKzor/d4MthsbU2ZkSr57ynBmW83CVe
aKPE3MoAaz3Ua+dmdbkH3LviXNaDPYdRAtLSceQnWR2pSP1mmrpQH5jQ+0eW
r6+OK0pWOYSbbRyZGrWfpi5SDVOSBhFwoByIVRDC4EHw8dkesC5gK6G6Dgrn
PHPdXODx/oZJQGJONzLwuOF+tnEL6mu81sQJFIcCwNRQGxQaZ24WCfMW7mZi
9ftTXunupOlXx0nfzXK7z5mvEN1HsCaSwxmAsLB/Wp2vxS2C8HKwjdjXd4AG
+tVWTxTtxm6Ol26N1xNLvBPru7HUHG7Hiw/Bns/F4M3rpKIzGonzOPf4nCse
YgJlH5hYMAhCONC8i/95Tx/bMWKlL2zui/wQ8XA3Y+nGDSJtuWmwrIQE0gmi
cje+S9RtwpjWteK5VZNWml5zekqNF52BcIj84vCs9beMt+rwob2+nyegP2Rl
6bvdxdBpT7oUOP36naq40CGRNPkFcTVGW/YnoVpbWmaU/+8vRS3JsMjtVeCG
3dhUrmCI0viIRTXg5hgN1mWm8OwhaoOtk0L2jjdM5xqhf8xI0G2AKvFHaEMC
BluV9dZkzY9YtXdfM6ZNv7B9bx619wwd06CV9HZNTyKiiIBF2/1VNG1d3hVt
hTMCaaEGtFsrAmKohD9vG9YaoBBdOUx/HZVoGG+5ssmccDv0PriE4MhqmS4/
EsVMPp1LlQ/NmZE+IEuY+E2ND985mpYUhT8980BvBS+ajZvMlRyVOSENiHrb
P3QSoPX4sUlCte3SMpDN9ZSV657tOURTSZHKzJYh/2gidan3z40JVHntQ3PG
gRS0uuSRjLHpnG4n0B9BNAuwcljdyYAZiv1w39DCD8wdjJD1Nj3V5moS3+Fc
+KqO1dEXJ70uA4JlvnilvBDx9+1jui/7If02k+y9zQ2xQVYTuer/UxDnqjv9
S3VYuBGBgZDLXnZHg+YVgfB/bl0HG3AUeq3oeyvKBeNSQNqJQgpHlZyhnir1
vOt2xPq9tLP/GmT8MPuFNClCmQzsiQesMKiFaaUCG8sOUZcbwxU6nuv2tQPX
oLGiZmpdEMBsUKegHFOxnlUtWjabDGCPoGOmb0Aoww0eeHuZThmfbQ5P2qlj
LVG23NbIlxw7pQPZR3IdMnQQoYlQP+3mQD0OeitEE3ocPjHgSQKa321aou6R
mQDwPYT5dXlS0Y8e1qR+3jMvuS5wqIz+cTyRmN+DezLHO5Xq93W9wIFR+QVV
kQ27KUw0zX5QetiOfaJ2w3ARZxthC83tMxQYs+y/M72bBobsnGBKfhoSsPBh
RtLdDusZWIUxjl1pgqj7J/SrloT3EmafsaTY4vOXTrHm6CuMkX0h56kce7ke
be5ZW9HxUSaMTS+WhlHeKgIyZN8ChUL0ci0l88L3OfW4AXBix7PAJYnF43w4
ekiQOrJMH7dU1b/twkUZNt/S1kGc+/bMuTEAm0qFgYFTg138FagGqJx6tQia
EN5I7ryBs+tIV0wFJdUGsSKVY24XfcBYANoDF6ZXz/ynZehZCQHtcTLTQ+Kk
nQ/NptKBZoIscObeODU6GD8c7uK1uOdl8H+sUUk65Kf8jtLKG9BoUM57TsuB
WPzJess2tu4k5hvmnuS9xCARmuZA+aFVrE9qfpCFRr9LauKvygdHLfIV5Ve2
FNCm/JYZC/De0PrZ2XtaoPJao3C2UsZrF3lev9gs1Mmk44F8j+MEc9M8ohcr
AvVtc2Aif0G0D04lOCaaxNjisOISpu35dIrKnUgsL/1M3AAye/WCyKoKon+X
hNwF2NAjW93MquPXwOUDRu28jKzS5zX9dMBPqV0jEVTy6CrqnQi7p/jCVJjs
z8gWX/p+kg05o5B0fuBVHyo8q42MURxhnukY8TbNuRat/VX8+RdX0lYIeD92
0xKjvwCYM6m+TAjIkWsdzAW55DTdX80pALK7ihTHxuBa2GnJYHMMOcO4nqHS
5bnN5dMNWbYJlcT+Nsad5V2dtUGafLSY+DqItf+q9SP8pXY2+BshXaF+67L7
MbXQBxJgm5YW9t1i6u/cjbEUitX4TWcsOIYNUaxP3R5TQx9IiBmO8sJBggSC
Itgbz2/ACaBZmvDakRemc/vVdixt8oQGLVS7nDArSYXk4YmFShcH2lnmTxH+
5zXPWn+PxS6o2gHzVDQ6omu++VJS5a9Xz0KrUAh+1pTepIsmrY65l1YXojFy
npw92SXD56ECx+5xaV9/BMciFmpdx+YX/HYBAwOqcl1sFQMmmEpcfzWJAdka
IPU+n2R2m1Sgh/E2KMjsVwGsGiAiw87vti4tZ8HdlS2oCA7AFa6WSo3RwDud
tYCuIYZvvzChJXks/ZdpIeM87wpNJtqUP7shodu1qXKopszujVRyPiXCKGe+
jHtnWueb/TYgsDpfcuYPntu+3c/uuQPtbcKqM/HPs6SKCYMOQhXu8zo7kbAk
qib+YBOhQtLwbefKsFDinkdPuzE+4fCGT1emJC7C1t4A8vQbUB/NSdCFCwuH
BZSItmrGAw6CiO4yL3iSrO3lVmtSI5kymxt6to5u78eEOTO2M0ZNLVEEllen
Z8iOHARhLhdqliMfiWaIztb7Fmp/k9q7I/AwQ0eECHwY3Nkw8MhfeyGhReEI
ou7k8PjIQS9rvT3dwb3/45D40iTDPVE3IjmtmsMZUusfKnQpLCjh+rvtsOKC
tMiWxGag9fy3AGiDoOmSqmEiKiwMINtFgPzHmqUwZKQcScF5BGpUOWz6Ag0u
1AyOgQzVMLuApIM+BaBdr5F+Jrpi0r5GcGOt1rmppMdMOI/WDy1k6hHXy86O
piz0RHWnj7IRtT3o/VQNIeprQKUuy7v9g4XGgL0L60PN3Vtf6QbUx6HGjckn
RvKWrkJOiOm5nhpGnU+EAZQqJfwc84hAliuIyIaXsqIaucAzfjanWG1sug0i
/NiKXcxv15sbLqLWNsYm+15jjOrBeJx3v7CyLfyW6HHhe5CYmXihrG2ZOi6V
pbbAWIPYTGTO7FkKyY3zQ/aij4waMWTDXWuMrk5FyFhIm9IZ+s0rlUB2jc3A
ksDci6APLm1jsnE8miB3Tl0UnaBq2fKSi0XnMxPghdfDaJjtD/cVya6Kqi0t
eLrQVYNFSXb9vE6phZJEvOWotLUS+VE0gAg1DROz1qwTYUG0jL/D0uCGu311
G+l9VpWMAAjR/mSru5fHFQb2ilG8H5/hViSkDEpbVbONVwVN5TcNLkzUaAra
jGCDBC4fXguOe/5/4qe3HGMi6bHg1ZJ3eLswO7LRgXdrnvyTpIiz5QNut3fR
c7YuzRo5vmwwvRB4dNg4b8tHyqXSWazA0zImlyDLa4YzCv910xCH5EYe6ksB
qPl9quOf1bhHY4nnH5s0eHqo35hYpbP8pOWu5FLvETl0tiJAkajK16ZMXGT9
AnL4UBUvgoFn9+OVfpKJlGlC9QqR11GRnI8rwRzbckZBlplcp7d85cFpXIjq
AU6WVOgFvCrlYmq2w1P2KyrY1nzLrygiT9LL6ROXPCHVVMdUoUQncKiGkLhI
Td2TR5u3AhhHvpZquzh0NWZUIQNn22gFvJUm+EoqjNoAtpHohO8JCbHkZ36h
kGj5cGVt5kpQhzhNII4clER8bOo4XQXHrA5QKlUQHcGICG07p2YGGgWxks0+
9UtA5AvD1OhpByEIL1CzjZWLa+ahsz98uJxdz9ZGG76ZJEo2VoXSBPBnNFjq
vrnLDRQh6ZldrDgyJ0GJY7POoYR8PV381BBKxItxNQcJC7ck2hKEOwF4DwGP
Yo7S3ZhH8sGCaqzA4+MCSkRwqBXj2Bf8ERuwMp1HB2QM71ACppGhOmiz6pcO
sFdTCxbGEfiHa3AXekFuWShYgyashoaomGi2+X8ommHStE0hh62AMsgwOgEQ
DlKB3zHq0S+xVi940WLnDSo8BbBtqVAt6hcoeNwKC/C7DWBilH0DRKwCB433
UwwP8dQxXgL+yPJEcFAEeaCM8p4g8Zo+Uj2jLEZr/LcAsN26Hn1FX9gUg+o4
flxpmOvGxyCoaJpQk1LeajA00xjqrqMyU95AYWcCNT5gkCfPz/TerRON6azv
LFFDw8Lzmbc96NJTvJbVVDLpIzji7/mhDDB8ua/fZlscC7wwh4Jze9P3zYLJ
vbNd3BEwbOOV0FIv2kCX0atTCfe9cuHASLEPwRtfYGSrK5k2O7o4XeNdAeA4
4sRcb8tMMKtSbEmEyWxTYPPrFmh+32jwE55lGh7Qq5NOW/AgtY25Cmskynw5
bCXK5BW+R1/XKUgNMo8ojcGZwZHePh8QqG9i2Qca3UUfp4qD7OpjasWZSNzT
izZlzYlVu+5H9eBC+fzZcj0bIuzPF5LFkrPpXxxGlXXqg7/Wp2bF0RY9Pi7D
eu8MsrgGG7mpK817uIhwpQThUL7RxRoRyhNJju+0ER0b3hPFG9Xf09WVGSLg
dk7mhJlb+dHCk0znQsmJWLspvT8viIxJDA0KYaxlS5Fso17CD4iDEuxFk5aM
nM9SqkFPcVQfx9QlQsgYyiKWdf0/6LnpzIp4f63WWyE2ojqThMfPm50lDtsV
Nztm2D+/1lw87El0rHCEYtyu3GC14uOVa5f9sikfFA+MsmNtPLNTObk8oZ8O
j27gnOsluoS4NXOmQQPk+guyp6O5gda9NAGPcBls3UanH3a5qErsAczyQz+9
iX2d/bFf/ZBr0EeubPMiZpJmMu4AxP5WIazuV4RV5Rb0I1P6rZhSV56bu3nA
HrrtdIB5KKnwIZyFoOIAQgZS+1/LB9yHn0jhkdfI7Qp7AR7GTYM6bpumExNO
5OZ4Xty1PMZBzVdLhSpIZdI9l9DUJIX68f55dbVbOv2N2UbOiGCCOvfWaLYY
OcHeaAk32v10yDsLOVO0SLqUQ+amHmx/Dit3i8BFZj5X4cGTDdZqnjmtBAAl
xslo8iNQO1GrerXyWuAVjFc7Qof4GTzmDTd0vKFapopyTgYRqOrA6cYTYzZB
pSbdujVtPYyudwV22bQ3aBmfUeQCXI1VSaxcUD2vGtdzagszhsXITUvT8k0i
qocpbzckEPIfmToIVioOyjmC6oDk5/4/RQn8fGHUbPZwb6hcKsu452nZxecD
rncFkAV4123ejp5uFzN9K4X9+ySilMe9sfPCi0L6iPZ6D/CI6FVOqsddDx8C
/1BISwsAMKOf2ozTR9wT2YO9bpbAJhPdpkLtJWDVvqyhVMlnJ+a25szRUbPp
AYGz/5Gd+W0AdtlTEjdYTrBHGkzhUIb7JE+cyVncrM/Sr8K6csy72TKU+V7V
8IqYpqwbk2YsGV0ocAww64m5DtMPBG/3Xwsxr82JCBDSVr9XTznqBDOsxL/L
6y2Y7+jNeWM6ap/j2EO1nC9otID0hPSby4hVff16bAca4Kkn+1Kadc+IbTvD
V3jc40IAzXvQXBvOV9LzFGGT8XIX+ftyqbZWp3CDSb9LK0K4YAf9yXdQnWVB
Ei0OS+J0N8tE+t28h/5hSTy5ZOZuoDTJQpIRXKHV4uySRTzahpBYkX/Wk9Ys
XDYdFw98H6+LDgYQRzOtH6Eg5VqXHQ+yJK/Lh2oErimDsFky0/dNeNN1TML6
EPr9+jZIYgXS5N7AC0ALAwXRHNH1yzVTclAPmwtKNOSEzeYMSMZv2XakaNxt
MzZE7eabeyqAPp+j28skVGZS7XjDAeCDa4GS1gAvwRULPioiXsbYWwfkkZEt
TVwFlIPT2xNLEiTdX7fKXjL73ycgCSROBVeYz28qbVujSFwgZU3M0Ez7/d9C
hmEgfR9gDkjLqBun0fDpqP8XtoT+p/E8uDcujlrJDPK5uHib2z1+Rx00keTh
avo1SnMh9ANUr9X2aCB/+0FTGTLzZLoAp/4g2y+0F7bnyDktSuGQcG0WN5q4
lYxIWVCcQjywTeNl6rcQx4cUsyqh/+bpsVymMprOgpivK2wEZjR00kOhGMcU
JgKMeP+trrpn5zSveTNi0gZl6LU2mw1o1uNGxZ+46QXfH5Jj+emH8q4c/RyE
87E/o8pAhibu7aPsKguiya7fhcasxUTPcuLIHJAqgF2Oiy7vd9YKKghr9zL9
ALGDcL+s8cpQZxv8FnZhskOkslQUAYZH5jkGe84IPHHkTY72VAhaGitadeOO
d1ZbH3mAZW/Ycvnaze33Eb6fbkqjKc0z7rn49A0OxngJPKH8mhUEdDrjnLn3
Q81CBrm9p19h2k6z+EH1qconZVThcEZgMF/PlC9bKkH7K7D/ZbAq20B3tASH
dmgMYiadwrRVWeGvSd07QQbqUd+rSZLm2W/lT20hOau6AR7w07pDGBPZ1kuI
7o1jTScYUnokP+vNUZ+/XDX2jiqmp9prQd3Mfcem7szEBeCdRGT6RSwQR+JH
IQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "OJXsOzX3SCOyhcBXS9yryN9cWQxQkhDHUr4mzQikLKNKnB6JkSYY9xNnmYkvVOJ5f3SnsxLM71tWjwpqmyTCVkTt4jikDmXDCnl6lQn2TVy78ivgbebFE/F7GUr3Z8AASPmtz4v12cD/Cz7nTJMTG81IGzEoV1S4KsV3MBcbB+1TqTshtjzQ4oMMPpNw9ltjOjjqx8CktvtqLiQWjnKfQh8i3R/5yQlzObBDq+VCqAO5tmii/GgZQgdZkoNIQB9QBMtN69TwSs/6Tim1pCeTcOhaLD5KgvnVSFXc7pZz4SZVlXRjwFg3A2R+GkBSeWr+myCfv8DJboPqBOqeanGvA7DyK3k9pJl29zuJT3ZoNJKto1WukC2Mp8GApBd9YqmolelTaAFYs0spNEcuth3cfC1Jrz0OX0D52hq7Nd39sjPBCTQPcsN2gQHkvyZPmPUZC3QEHCcdcDo1r4Fg6kpogy8IoaQnC9rHK2Z/RdBt5oAlTGm6dlNrJIoyT5UJqV6CD0YMGS7wpWckJAwYHCQw6SpHudSL4gT7oPbwspwga2r3hhcG8H5NyXHiUvI1tRaeNKD46ve81vuOco6WlWsieCZ+bO6yWYANYt6wwa3a3TaaIGnbVeMI0D4sFeMf9shzTNJ3Fhu6C14DBMa+0TFppc3GAHajKfMW5FcYr/4y+W48xv8OCKf3GQ2CWrIbQsRBf88HrAfrhOLm8drfMnZDYDlOTs6SlAPq0K8sdAT3MtuQt8c740/0TfoWBtdNzyyoBljnH3YYHqgTBT+G6mzoaeokj5A/YHkCZtbTFPc78IuWXCeXlPX+qkNC9m0Mq/jlOnefepmBuHrBZcxdh69QljvAo2Cpd5NApkxtGuP2itG98c/G/GumQUPxGl1Hdi2msaYvAQ+8v6ktrl/JImNwSkTbiUHytk2Z1pDgC3FsW22+zRHZhDs/puYDpoSTILlJD4MudzL3f4l2sVlamDbV0GDoaNJ/xcrETP76Y8lBFo1mI5ZaCFNfsrTLIOWrLZA0"
`endif