// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QcxfY5N7HH7+erCUm9xzttYPKWvierHH2ULDihHAJn2WCCjRYVN8iJqjHD77
0ProuMy5+a4gN/4oP0YY3ykJ82otEIY5vxCUo/EiI/D8G9q+edne1mBIVzTw
dgX6h80QL32MfCMf7rCTwxSCV+gICnvf4jGTynzFCT0mTIUFLyyaWGNBhZ34
BggSrsXd7Y+uGyRZQvmIkTmlk52mAsrzX40d8RdVAXeGSJbtkIvkL97AIYPg
Zy2aKc+muo0ROzdzPUZXyQJILmS/5ZyPxK83J5FEik5QA4rB4HIDL2IFcXMU
HOsOvaPEMIeWu0Z7w/p7SSIbih9DJMATQm+zLLMW0A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
C74Fr5FCLMJndRxI+hTL9YZc1oRDke6iF3z9n82UpfEs9VGt9pR8q52gnlP6
VJ57x4AEKRfn/YVn35mkP9pIlCIKGnYBhz24/Gmw/uIDXowJZItkZrfl7cV8
VPvkvdT4VM5JWxs7lKJkgI8FY5FgiL9dMQ2S2Yj5b331ncsU/BY3LEkwfdje
9U00Q0ZSTdeEAKm+8fdklKCwdJVMdkRyi3zD/2nzsfNDzm45WqER7n9ZMMto
xrOz+9vBW6zw6laMlEF8ylBol+2XYifWguivP9cu6peWTfOnqdq341OHM+Ms
EERaAhKJEHEMtdiVyT8umWmW3YBH6LPGbCIKWurnYg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aoVgxyk6DeEBBrHFU5LirknPlKBkN5cbU5dsAKPsAv3rQ+Z2LNALmCawcM1u
eaUW4EJ0t02PbL0MB53+TjFiaTiAae9n6CY4BQA6VFoI6Bh9K5atjqqG/HB8
ayTRnW/mKOQfwokiQDVZRi1Bj74CbAOoC39QwXMe9fyrUpMp5DM3UDGGWNPY
DQQeKL9UrzWGVBfsxE4+PGihR+0V5+iETn0ENUH6PqCcFy6Rfw66WQ36qedl
yZmxeFw1DFEHFAjm4mFWW8Oc74WriFNI+OaqXoiYTUocrDxi+A5lgpowD00W
hxom+3kcdMOSYP3ZeJQ4WLRpQsC3byRrFKcw4oxarg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MO6NbrZGIHAIL9XsPlV6twOlK0YBlFQ8a16qGNzCVyASs3ygZETZ/bCpxTXI
uFJ26ADt+GLyiHUS9pST8lftk/IZ/dFAuDz/bIk1LvvvMhQy/g7gTubI768E
9Dc/5zZ+gxrhq+q77pGAb857Hro/EBNpgUBsuQTwaUpbJeYFBM8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
UU3EYoGLupnEQMkU8MYYltCFL0YOj5hQqN3c5CSteZ7VyoHRqfvRF0r7QKUk
CR9sB05Fm4UTKSlA79svIdZIpzjYw9SGoOh9oWR86WBh0lU1dQ8rDc06a9rE
oqu9H7HUeN1oc8FWy0nKYMGLOI67Gr9VcSGKmJhr5d3YJrKH0Y5yMbTtkqVE
kH9/TeEx0iUCKuPnjfAzHiVyfEKIHCEMlRI+SXQUYLkzh6lv/GHgn88NXruE
r+QNf7t+DVKLDOgH6fcRQ31n45yoqVvdJG9jBwSVM93pwJ2Pk5l99fi2e3ZA
OSlwbsZqd0g5Cn97aqQQ0hlpip4ezBnpq+pPeEOLE6HecpuKNeS6OKAL05iC
phgGPyozBAqvZjdO1RM6k5UtejlXYzNRd/+TlrfDP9vRKso+h/HyS2VAM3b1
Fx5uDMWaNDj5RYpgjhw0eqDTMPaCT5gFEYBApESaNDCAy7ZUsvM7/30xm+Ex
NThgbBc0p65pnZ5xj1cscINAVSdiC0qy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FK0QVMYoMyxDNlCDfAGMN1G15WoLmJ2U/C6urUyPT7Kf6GtdzIt7aKKo5IAV
3qUyZREjPBAWw6ioFk+jhp8M3A5aJsLcjiI+LmJzkF3Q0TlGPqLzgI2vN2tM
jpHo4+ECfE5QsrgKXQGPC/6OwDfQ3G8/1xvzEDY7sAD1AdfbVqo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qT+wNdu675l3S/lohqwr05U6rSppeq/gPo+Fw55Co9FM8zkgbZL2dxCegYdV
W9tbSYk3PhjKBpcRiWKj2jvaBccSftLEvPM6pVcZNzoC9S4TefXoMyS5SgN3
nEmPnpQ6OsXUQ+FKJ8LaqISAx8JDtuWZHMBHjUdMlAQ82dplG+k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11168)
`pragma protect data_block
AnxBnaM9EU3w+Ui0zvEZUWZVsCnEX2xsS1D9rW7Ww2/fFs/pER9Y17TrhgrC
h7m912uoYAitwySarlpFjozxd0AmQUYpNQK2DN5Q/dVni/3iB+R2JFGnJ+f5
leiURAevKiMbI3d5xeOuF/WnzTWOzGccx6tIV6B6JfGy7d7HSSG93LigHtxT
VvPENyVIcaqDuEhbva3Ajl18kA3xJRcr+glSNaO6rBFiv9i/4opPga3ykJ3V
61VXZ6CjIcOK45y8mTPQj0IrK/aSr4AiWRlcQ+XBFvnvw0ibm20796mpCZfZ
szagDZuqnYVgtTxXL00AB8GYyr/LGdRGOIH4kMZFUB+twSWbhbq3J5alydSx
v0IPkBjiXIDdTXH9vG24HElO1MUAbBXnL50sApgsKPO34WAb1RDY5dvIxznL
xyuymqnPG1NHEtqYYjavnBqpRhFcBDuJWXYImj23I8ClTxS6Ccucl4NZQrG7
37/C9wWG93kS/NsPjEafvyLaEFIdoCHxFNv6noOWbjngf8w589BYMFVaDdzr
QOz7bcyzYOcBpBBfUhHo6h8mrCjkk2LvvIpGmS8cmf1AA2wnGvuKH+vwVdSq
xpGUuhSz7s23ExMC5bUTR8dDIGeUWg4O2h5zlpdx94wBgqonLGsQfylGYhqg
5JGjrYGJG2deIPiSMAjKRaw9KBKAvmHbIqykTizXXGGi+HzJhlbhbRFpUyAk
ojAHFwSR1VSI0kslcgqCibcZ0N8/r9fe0y+NjLsTzx88h/yA0Oa4tdO5c1Ch
UtGgjWAwU1wG1lOo6/9gonDIDxef/6B5A5vLinkXG2snVUO/dKC+ZuOIp6/g
ycJKXQxB8S9oiFFoxMifMYF9X7S1xHVbIa/my9CF8z9bA1BxlrUPBDLQ28On
eEUpHLzTesAlvEW/NJAeLqXxSO98TkeHVGUjvqgdqeBomlnpexgkQ+Vc3Y/p
VM2Vu5O5iekbykJnh6McfoO1mHAUeoAfez7upk1EbcB6WHPrulOR/ASjdE1a
jt1PH4S1MLc6varO5k4vm33kJk0q8DLDH7G7GDcXvt3yL2rOFTnbQsbbCrop
NX5Ahp8XRCaUUfB+ibbBFBUV39D7Z7I954C5fXmvuQ5ROccc70voMeiNRrC1
OteEw1kadS2E8hAoTvRxYU80y5cDTc0OT1uPxJCacU0mpXNYGt5iSDIswvtr
FaDxiKgiaDVU9735HZjw0F/0QVg00XttcuAaR910e1EkLLgIZgpg7q32D9LI
YzhEcQQulsbFAo8O1OrilRPQpULk6KdpK92B51UGjYHiJMDJsaSKHTDdBRVS
GkIdVPcOnSTsdYEUs4RH+qoo8Fwacv6ChtKEQn7HchuqDyl9B88eG2szxzK/
luFZtDoBCgtF7JB5vW92obj37GVRLM1yaX+edMFAAGkowWUQts5ehvDx3b0r
B88E1fSQTd1+C+d2fnkjfUJ6O6ZSwwQhKgGgdqGwIzWP1KGG4NEsNm/K74Bf
rwBgTn6AS17L4/LIcDvl0izHGXQkamXPdV+ufMVCWRPFP+An5EwPeCY4HC9p
oDycFSYOZZ91ytbvB9TKyiBRw2ijvrU4lLvtzK9j4v1+pEQnxHhqA9i+Nken
hffHk/tcPmUtMo92XmVVCXrbjIx5jg5o8x6GXl397w3E2u44v+qkbOPXlL5D
ScubTwtCOsMKOpZ4Helhv45BmcdqvgdYJ98oXaRmL2XhFiGW4FTbNg+syHBO
Kyy+zv0ke1m7IMAkgjiX3dx0vwbpSU2pTcu+PIZaXziSTyoR4TGsLTFrTv2c
23HQ4DZvf8mA3jiNRLu8PVKfZm+Di4mOaHrbCWvBm/l7EWzQmMxWZt1ooWG2
Q2RszLHWTaJASeJSkEcl7MK2m38VmcVnAmCWwc9bF66fDWryq0MqishI5rMC
Ry5GUwh9QUig075SdRFNKTuSqorLW11BytpMMFQ0ZX36suDsKkmHiTQXzpC2
MGNqM6jyafLKzP9nMs23qEmcjZW9lSAwZUwcl0aD60QWE90kpC1GJTcceG+u
8+QpIXBNbCKLXgDekhGhSiQemOrXcSUC526p9WGWuOwk+Y+WP0Hj9mAJHRf6
5GBeAFRY+E5465KlibeuIJnJUvUFSwtdUU5PuCsHw4dPEyQBX/T2Z/zrB1oM
Q4M7ANBqo94ERgHIgb1XaQN9TiGMBKJ13HgzAL+cO73AHFlx5n4nAiFhcWVo
m8dNmOPTBvec/XWNTxpYo73iApHz+TwbUoiPw+piH4XboFmJhyoT/uqIAfYk
/HQ/NDkkrzMLch7tZohkhBanyiho7R0XNRHVDvILF5q1bGCZlmTfeYypTp1q
gM9UxjzOF+rhQRtSGxdtMGQjy4nrFeAyv20s2M5T5/8QAOQXyKEtCWvM9crC
3w2EihK/t9tgqcvZVE7vJ8WAoR/S5+fd3B+CCYqQSnIm3tcLB1t0G1WMh+qH
2y5duIccQ2EIhd7wMkRKRZIPeTSrYa7SHyndcv9rlHCzyAxuxWwF0PE8sgz2
1jqWrGMOgE109alm14YmsWkb8UlnkalGE6gB6hULRQSkdj/afkNKQ4OFed8T
nUtHjSNAHgW9TLCegYhsJO8iVOG2DCezhrLZ7yD4+BpUuCG6Zs7Ej1LUsjRD
r72WPOKoaxBmT7Ms+9RAY6EMtBSl6xij/B8TnfzRXvEQwDBev3fZhGzxt93b
JFSKKOmHUmuhJauid7t+I81YsprM8V5whSLVmTwWM14k9iN5nstSEpK0Fll1
8+30rWBMmc/d4YhWcqbhnxytmQ/UOV+ONfUXnffGEtorotUG5pdgztMbjWVp
Fb9MRuH0Xy9SOAS1V92ScGIe30k3TyZyOoOzzKESj7fLfkvEpHISGP/R3xBM
5RAgzSw5NW951LTmiv4gyFxHutvoiIT9YVEMbX2FfUUXLPq3Jzy0sVMV1o0a
wwA5SQJR+y3BczBJSGQACAmU1g2LjfHvezGY5nItTSTEntwGovOSc65Nj6HF
ArrNxh4nRpIuz/gdaE8m4/CT4FgpI9l3sZplTM6OW4sv4eI1MUqheueSuXLM
BiQpD7i8f9zd0S2hVKsx+VoVhyPnbY9SXBM2VqkCA5cKcsr1d9oUJZV4gDDL
n4Xk97OnRlblDCsgmKal688Q4uuPZOIVfEb5TlCQxC5Ikt9IeatjmSfjYvqh
dh94Ma2Ume0fEGx0ojvzbKXfBUCOkoiz95rYK7QNg/ltXLGa3vmtyn7NebbU
sttZ0IP/aU/NwMF4DNG+EtrxsbTkRLtr6+ONHhukqjL+i3Y3Zr55wMV07EVe
I2bC+SA40XWnEdiRBqGNyxlQHUCR7S5sskn/Gi/KF0hil8CAWxD1G4fTkH/+
HfKD+DkmTFY+t5V2yxmOI+edLSvuQvsgrwbV1I6fCylAoez4/s2n+6G3Z/ot
jAC9oXlpTZXHqpaLDoGxUQ5uwBdiOZL37qzMu3NN5149Z+OugJjXJZXZzuko
EvUTNtf/RxlrZsL7BvtAOEtBBXGT1aMtEoynj031LDVg+BGyEktfSemn/pnl
CRNrCpSQ/RCiNdaYWn+WeSaFZo7/onSDeETgGPM1xJYRNw9rT1qBBFh2Nvnt
QE8zWAIEfi+EwYiS+tV3owHm/4rnhJ8EHTjpdoC0XRDlcZrJ3vGDxPmOfLMj
lSGZzNjbCq+7p/wNtlaeJE/cSK11XN7bPivcXRDUCBLehf9tXkGrBkBdD5Th
vcNt7zS9HLd7tBIOgtxSHWzxBLqVntWEKCcwYGrN5iKePvzebsjOzuCtd9I9
7cbR887ooPBBAI945zDjqiVu0eM7a1IcqrtWxEHFzTJUQJb6XCKgzAyirA/q
D8LAW8XiDeQY7fTBN2FI1GYHtWu+dvfaEqZSYwyDsttG89pDoDxIrVDCPNaV
0S+9FeatsWCPCFCQjzQPbGdPoi7xaQ8NsS5C4xa0oTtcqYc4pvFAaKywjpQC
PVYqemo5B8BWq7/PNvQOazDgtIxDt+tB6qZY+hsHZ5I1uLJRk4xN9GZiS5fW
fO7r23rjvgUoK74O22vQPT8x9UUZpf7A6RIGf5K2Pa70ATOfmYHKciBdgVNA
+mD5kb20Ep1xD0aaaNCn7INdcb8M04JhbWkYUQtbQNl2Jq+BYjsUY5MhF5XK
OWq+tx9SCyuiFzsizkD0V2dGyjwIrkM19VdGtyFG/NaOAtZ0daPkeVbsXr4n
CWp2E1a0l3czGOM8xX3OhUzURTmrLSqHHVUGDBY7G7Grti9FYThYBU4zfUUk
R18s51o48effA2pBV5Q7B0Mp31Bn5dy8RsYXDfMQOsar9gFSSAfADeEGCXbN
gnKJbhG3DwjFBSvRfgTlXc4wdog6NQr+Qcph2UzJrKuFvUhsmNYs3vY9uxKb
ieNJPRW4KzRJDXp7CLa6+oijA4qlKaV6FlAgW9qaQZ3Ms5ZHyXqs03vbnTj5
6OKxMQ8kupberYHHD9UYGaKAQs1ZanZJhZHxLJ/IYfAHO/ni15w++GcyAzOG
Q8yAVqwUh++fkiJtchltSR75GP4RtkaVMnlvD35B2wT0K4Cyw700wITMf2/t
qrEFjjSs475x6bPP02STqPLxf+ff7fJcz/3Gs9SplomKTDvyuexyvh3zMUNW
I+5NGYyxGKxa003DTjnczLBXZNBRBDcnQD0JiRZNhD9ru+cn5qm7q9uyjEAH
rGQKr00qhOyXYmmgrSp413kxZPf/zMlHB/jOV/kT3KyocLU6LayMrlrnhCD8
G5AoYrU0BMOhb1tcSTCi+oAKamu82fcOtJ+wD+lpOreAUKcwzm7n2ViykLNR
Iu+oGshRanTumZBVSAlsQ4nQOZwxTvb5JqzGeatpPC0gnyDBwTo34yqMVamU
kFNKmN1OaBL7YEwCuD3a6vDiJPQnUobHfSKlZ3ou2xO+ZANxNYUb0yWsTOGB
3TUF9IScoA/YQg1qRvHHqlNcdTTwGgMbCz1q4dDfA+oAbHCgUM/gv5L1xHMB
rr3a3KEF/YFwxLdSdzHfd53uj32YOoFEUydDO2vdfnRpgC8RAk3S6YL18XQk
+b/zj49WR0Xl6WCRljOy0wOAi78c0aQd+vsewbciYRwF3XD7HbScTKh8nNtc
fJzSi4X3TaFuZ/ZDqY50BfCl5KudBHDPX0oxyWZaZ8pJ/FpXi3BqrxDORWjh
HR1lGVJnVaKTB6W7XLxIymbu9rsMnYnCJiWopueoz+PhwRQiL/xqK8j4QBvJ
6tNp+zbZ6WNrw/+lKd6MGNjxkIJSd5ZDiIhZYi04DExMgRpCx8gYnarS5P6R
jxQ7uOrOKH5r8B3NUrMApYHeGN4h5J6ps53BAtZwh98DuyBlwKO5vQzKiczq
9NuQANcJlpSPVdQGjEC1EZwAplvFDm5Q8n9AjicZucoMjS8gpYbkcCe63EjY
NiJXGe+1TY7Gy21MSaLtHPSDj7ZZyUykjgY35ixnBOJaJ7mvRrUqR1Y6CJUD
dnVizsF5u/AWyp46x9mO8yJ88WQb0KFIhxeUHR39f1miRjLcLyx82h4hTR7I
MqseRpZeJLEJEHYZXipjaeB6BON2KFltOsJRlLZO1mGWQ495klwr8Wk9GOy+
h9afoVDFRqeR1aAppYfIV4VjGCdqEAphT0zIy6dekCiFcXkzJtfXv/Ofn536
4tZQR9SiD6yBdgOez4jBSRNvjHcXl6FGB9XEeA+plKsrEePgrI0q/b9PuA6l
a1BRLUwr1P9BApeqbupz48/xN6QdS5g1RaQF7panzEWY1R7b1EBZjOWFZKsi
nmuT+RlUi0u4fc1t92749345ZscaJ92BpRffjkX0G0UBHC5TADVUgKBX5lbk
chZxDQdeec+PBW1Bi1lQEvtN+f7MAgNL4LOVD6uj1mY0lrxWcUsdLDCAN1Cs
g65DWNo5Yo7vYJkyt0gifGMCk0hnrDt/B8Ny6wmB+6KCPIr3W3L7+KP4P7fs
Lgi5MfdzwlmAosSvifYGU9uukx+f4w8TLqG1YYhsMuZJFALCYC8zfxnG5VEm
Gd3OvMG3ZllBzibpVq8Jj287MKy++/cSJei2RR1MdiHApZXsb8aaiwAe5QfM
zoBmKAqbzCSbkaxAFORUHZnrwEeN1+2VDk0y6VTQRE5O3tFgDwFUpr7xc8fl
XrtVxhPFrAJ5cUPtMc/utXKIzkNFm0fOCemELZOMZr4OM5Pvq44Ic6rX8YtC
8Bg/8OM2fzTpXE5gIrIySd9Z+D2lC790dCstntPOuMiyN6KvqmPjOP4VVktc
fcbUCNjd6ZYByQI4OW9x7enuBA1mAcjTrJJ/il4Q5t6F2oxOFolw1JjXfke4
1CUl9GFtALzC2ThLwGYQFnQrs94FQNFrTJ1Ia1vOzP5sj1PXwcv91MfWm9Ou
hrlpb+10z1CR8j0xSzSyb23dhg2k8hBiLiITQWnqzvlHJwJy+rB/D289PqvB
FshUU5Tfm6uZGVfJIrbKo3nKN6rvReWMr8s9VZ5AD5cO5iuHqfGTAh4kTb7M
HeVA5zzwGxyCY2lgkU+hv8AoDJAANQafOWK04ZbQD5zfGOHHcxPEPCNcpcTy
5xm9Q3Eyu5hOyWysJ5numgpV4MAapVCHVXE3Ifh0xB+vZoPcLwz8SIR0Py9y
tpLN+dIheyoRe+89PI/iZHH6SVJ3cZ1URd+HtrBuWLzI9K4b0CX5BgFaO4xj
yuV7Jw0knVIPtxFNvBTjffoWRFUP3Nsvoy7ox0Ka5R4iKM45KPHoa/ZCDaVN
g7ReMzCpVxntD4Oa28QuDxzcYrpscW1koXs0U8vzna/UgfD2JcmOAUXh7fxv
iDshWx4otpsSiNTOukVRgy1AQktVAIEZg2QoyIq3YCGtXOcMKZwkw3KR2Mga
V63atTKZYam8735IjomuWyjy/v1d8LL20xN4Dg8CTL27yQysperaDQ4yVL6+
A7bP04Tv7RXSl3TabZqg1Tzo5wyknPXYFWlNXsDCtjqBHxaM94EDBHz6VRgA
0/blL76IEiAoTZubJ/FJPjT2m6Pa2HC99QSZCaKFLlXoUCQi/JObMDGn2rlB
GwKliNpA73d4dbGLHutSiK1xQCjKzR/eSaPLDD2jH7gQ2EfLOh7R01ujnPAh
3qOumBK9tc5S70ZYZAVU+UfICq6Nt6BTBgFyNXZj4gCIvFmgjgoDryQ1zW6G
SspAjOYsD1qFe5noJJTnHl5ZcbmWn/3oKkrtpQDs/IN8avu3axTKRogymXMr
X4F7nDQyTYOeySRc1l0gWKMUNeKznubnkfkv5/3DiQkwdvw8qJAHxL/q87Fr
OOclisKEM55VQT0zhxe9RQXhUaL780/A7F3hR2zS1VwkUDDUiDzM+ij1SOik
eA60KBGtFbOM7cdB6W7LIHz0ry0ZcM+l2wAHbF8yG51ueDvEXfNm4k7ewpbv
TIl29dUFg5LhpZVOIHxplsmyavfNFTOQpJR4uVImBFLNC3G8FcuHypYvK1dA
Tn32ZN84+cFAeiuCoiRXPaiVSDPNb1Sbn+pPAKu92FmRhD5nqOdvCcvFkakK
Lu3fSoLe15t+MHa4XfoY20kdqVipgv/LN0GPknbfO2px0t2ksmjp8u74LfeQ
TplzTg/1ld6nwC725sh03sMW83xYgYzIiU+znFmf68zcQCTQPC81byJ7zIcU
BCpc7WRyLa1HTUTfjKSRYWDcwYFZU4wWzsNE8wvluFxtHd2XqpfZRyXPLyYF
ojhIQ5vm5Ss90WyM0rEvDpOXYX/DYXIvWlQ/B5KKQ7uFZOmSb6KQQcyhqUlU
UEAfYcyrdCWUl7ACrOgRyML1Innw0OWC4j6nMV2lTaZuCRjauqCgbdmTgJnm
e7wcJpUtsBs/Iy+G/s55og73hU2I08YWRdaGFYjjB9OYmAjNvsoyg6Gr4nVa
ktrZLJ/FbAOJHjskKFHP5Tg457op337VcCWooUDj73tqPIsvxDvgdDlgfzLd
iF+ZRJPxj9bCshXrXL91GITqyy7dt1/KP+AkSvvL9Uc1hWcDDA0q8tl+xrwN
8yreJDW1+nqvFXwUnPd2NFWRiASqJjMDUL32EoqWfbYWlibOIV4TfDmp+xlA
4A3QD2/6U8w4XqeqYgYkTFfHm6/iEq/0VzESFSf+5t+SSZxQyH6hUiw536Di
AD6X/SD1CadHc9F6+Qm8y5/RugvUn+P/K7fSbov57IOVF9/zzZZySz1ZqZ/M
xIZal4iar4D0kJxvf7L2Po4xEC28RrmSufvJoj3tIvr6laXHkzQiVjhzXjay
wY7Yp70LRIzhJOyr7H+KDbz03A3gIa0E8G9lOzorSFciunX9lR2VfiUBLhNz
NImrYAeWUxoAeu97i2OLJgAUlfCsm+URFg94xDrB2D2W5KlofYOahCCiPlHX
kwWhFj2nwcgNw1PsadLFy2I/MRoTpyyxU2e9Hy9w1J9Y8Qn+Lu9eJUu+CDC5
lkJ/aWBFSbM4et6VI6Vw6HPFE7ifEmQ5N7rbzlz9DHUZ7xTC1EzKsjKbKZL3
LKt3B3JB2ySkfsx4ipuE4qpMxxeSPbe/92ryvt5mIUzd1EMM6xZG/H2U0E1a
8RuuV7XQqRPfUsJBcwJWKDeqT7f2NJZWagV5JtxWnxWzKMUl56vdeXkzXIi4
T8AB65fIVKD/ZFkhcO1WQEk5Mqedow+I6+D3kI1Powyqo5HUJVaTdao1+GJ3
xVGLhqUDfyXkb/tazevc4Pd8DIOcVCMoNpdNjSuY7IKPiwFXtAN6hdEe1rsJ
4s1DFM98nOvBLvJmllCzl3ww/q4tP5OdTsyW3rWQkEwSQCxiHMYkEE2pZGlf
tp6wiOJNuUyG/qNPiCh0mZvNlOhXLoSyIgzw9EIcq/uoUH5SN7gB0gKHTHey
0018d2zLnwoPR+vK5nz3VcwyBcPYvwlqDTUmypuTzuXp6x18GPAGEZI7OsM9
YiLGOQ4A8ztZxGxm4/wTaRcwqcxb+Wu1DzPElDpTBD617DtambnqW2ulz3ZF
EJHa1ssb6MguRsfHi09hgSqDlXdRIc5nrA13Yilp2yWp9RZxuS8StfB0RJv6
WLKSD+7r2wCMhN/OjlHwmeas2BfrsY9T6efmsCLwUzSGGgU1qOpMVWLwpaCY
9hlW6m5m9UzOXssnaFua7Q9pQSWBZ/7/06W9crWLXgg3yMMiRWYHZJMrhUD5
7fIBPzKyQxiD59mUw+U29o+gUNXVzANAIlN+q3BYK0fJo/JiS3EDRb9UqvKx
Y9kGdC/FK2GfStPBoCvuryM/UQWoL9DXhD4jWhz0Dh3fUXeeQ/vIizPMQXNA
pSQ334fhPlTkafPvec8IuxbVc5iyoWkGCbtQSM3CYzNDoVZ8u6qR6Vc/DSoY
jN7fpgbk45KEm6OA1uPnR26dFnHIhry602MrYmVgufN0apZjYkIzPhtJYgkR
L1brDOZUJ44tRGIfkEQ8os3+Ru9szV8IbASbhCfiS/GqusL42ACpKUBwnSMv
XNIhe/KIp2Qx3eFNIIiJWJ9yt6V9Ias4ra8g9oufUSLgeiR91m7rMaAlxJ0S
UPQb+TKG+uq00lR6DWHyHWn2mqNU1nYtFvWMucILuu88xXQ78x/rI61DAoOR
ZbiuiaFfskmhocGI0GOh3+lTWaYoNR4Y/K6TclPEFI65BsRf5XarfVfTSpNM
cYGZ7gwdyCZdSwt8iJunzdQHEMppcuJ4Endp1fSOJYvrqBVGt1WerVgieFo5
DJ8377Kg0pQGOFxLmKqku1y4zGQBcv+c7SNXLm/3XHzYYvWPfsXvVIlxohR6
AvgcP2RiRcjxaZaXaSmbI47J80NSKtsfyfXktkdVq10qXCFPAIpes7x0mcH8
q4PTr34X0/WYxKYJxxTbL8S8FOf7m0ZtGxzTuwDB8couEDueKLmS3LWjlbCP
B3g4d6Nh4BOeRCOX17C03IOQAKidC2Mf7nIZui5Nwi08FwcVRliFr/JO4gyl
Qt5CHP8SE1BHmgm2zw3lz397fpX55qTAbxDwgWCEKwOtX/UKkGGirAQsPoI6
d9On6vpxC+VC5MBu5bs/Q/bcs21vbi3/LYCd55D6on6PoJPFlG4xobIm7BsG
HHeTU7g1MBZY04bf9HevHlx79ysWEL2C4nlWgjZUqZKiW+tllNSnagS57tif
9lbhwjAOcEOrWYb6HwOKCONueucxNACCSCDIqv5DS8cpt7N5KFysCkrkmvGo
zyGVAdueB27GP6BQhHF5+kJPp9CaW2NrNP4n6nudqkDiIQ6F2di3swgpMArO
M0rhAIy1SNWneKPXKBm5O7Oq+2NNXosXw5gAdcsQAEYD5fIQHfA/p77KB4Tk
IH43BYIonx7kuWt3Wi8L19xe6j9xfJBGHwnLDnLEYOBR3PhHEBenniH6DSH7
bbePjWrMevg8wlfWUqsAi6lc9jm0qknjNYu05gFy+uafL6PdqAgZfMjuVesU
TjMOQ2ovuzrgTnQ88nVqvMF2drOGMuASoqm4wE89SmwTDg9zt8kOe7KBP4Iz
tsr3szB92QAMZyK+xrkwoTaZp4NYzIWFIX5grbOCjyZ5/cCFoWCdwddSQa66
RlY4t2Zw37ylYxSLkbsj8WIDFZwB4iLsF/Px3klZmoD1YjB2DZkU+v/SGUAG
f2T/aJFE3GwdhlVyfrDeMUObHgN3jYV8QhYFtIXm/gmMfCktptcht7rPZgtq
4Jc5Tk42iQ6877FVnQdW2k2icUVw9eDf7SmIb7kowxyORwwr4Cr6BoDXdo3j
hJWweFY4xPytZ7OqcjGQAaosfg4O5/Dy5X6xdSx7AAMJVGKFVhbCh5x43mgp
mwCmI1YTlOTupjBuYCs27HgTFpMxAFibrKiyc70gnWEzhZE2Y/jA2+43EtAM
xytwpY0S9gd9l2K1hDKymFyyovhVHVUBYPAVRYrYHB53+KsPN0dbp0iGvAGv
aj+rN3akPf6t4u5GVTMu46dGp16pF/aXuIlZnc6oqwATyg2kL5eJvqbK8sjj
q8tE2k5TSvwgk3s+K7g2Mo3USBMUAZ14W5g/zjQoQt+/kcOorpgYyGDUemsq
jpkULWuOJUn2/zeW3dn1MvZgyS5xRMtVnOUlrmb2vl+8AH2EQL6DXenQA1Hn
wFK8bROqcG5mfGxGeLgJdOJcXvPcU/01dujSHg0CgJrGmEfZl0ub5nV7PmAx
AG4ZbQpm3XPEf3SJdTdSeQbbLTChC3nUYgC+BpVwr8roDRVvMOXnB6Ym/12e
7+LrbAhPdJapdFfg8uQrFKIoqmjI0PcdKlw+XD4ZqKy2bjoVdUi71Hj9gi7N
0djW0MmkwhKX5W2OAZvA0LwYSG9ri2T5q4137bg/wHyoN5r/FBsdynzvBvZY
gMdspiu7QvLD+JQZerbIPDd+z0V1ku857caPBEdTvYImBiG5IjJ0yPcI/+Qc
+4Fu7Fal7V5wOrgowpuAnd2dNjUDFRuyIIimM2s6QGce2Hpd4+6fiq27VsLo
eJuLsgxJICa/+rgZKuxAsT2DBbR3VrUBKkwqo5LCIFqzErGkpAkMgLYG/CAM
jff3YtwETfPxyjHhPu59b1dZ9ML4mZJ8QLFB4lPA7wfPyZzkeUsVx905srOs
xkNANmGIMyyJ4Be6LcXcMAvMCJ0yrmvywQXMRHTfyZdK/NFI0Q4fH42jjnIS
PV5xb9IL5owtdSbbx2o8TF3PCRfrKN2ZvdxyzgXIIYjKvZbjjYV7maYvGjUz
+xLftMmJgTp3LaHxrBfW2qIpSkbAO2cQ9zKYrExY9kKHlGI1BhfyBhQ6kuat
3zApazcjANM8l+sg8XJAdc5R+jLMDiT+RpCxie64oH5uPpV6gL++Qt/VodN+
/KhoaQ9Nd3JgBNhNxw0M+0LSuov0opgANDBdRGwxSGZMHGT+9eNAySVQQ8Lv
if1UWN7NvUiddlA8i9vrH7dSXnQ3E84pDdodBEHmEddeVLTNnhlUS6LRy16V
l4zFgsNRkASDvqAPbI9v280LRBRo9lRMXuq4jcKF2IYLG9NSWblsPNXAuOKr
s6IvAsNOdAxLb/6rw6oE4/BmK/EMNRiFUTq6jAfzfzVqMuqHhOlNF2TCRoQr
k9UtcZCb+HB3F3tAWyyct5UUBdYliRgrPJbRSbXSOJN+rTkqHWPLGv/pTwWE
5ASMobv57+k8VcjvklCp43JbrJM0KWFkDw79PEOj1JKY09Ih/h06iPNm3vdl
uL74EuFhIzkH36XnqJyv9CseFrS51TkCZTqWAQGv6AXzAbH9BcqmtKcXcaVG
FaVguNeilGA/lPq0uBKSu0o8B/GmPSz2vv3D95BmRP3RMGbv+NJUoMgXzQbL
CrE/a4oOgUR7QmCXRSHB0YtmoSoah35x8Dgql2IhjoyG/IC09DuizWIJG4n8
84AuuHV4y1421HrcnIT0ihwTpKThLt1d3COJ/Q08xXHcXPm3YROXryz182dI
b7aMXVQ9FajGa+6GgZmSCoNKKoz16oDCWltYYmcnRD/cIKpHnRiFm2DuWijT
vskT+/G8e/GRES8BbhgEGNiwuETVErpydIaZw1E++MJLarIQ00QEd+8AcR1w
Gux34BOpfFzzagJlIiwHJN3lpnuvLjlGOZ24oiA8zuaqQVS7Y/2dPtsxfBLw
Wz7Zp7c/uKcQK5XmMi3o6iBhtGXHSwu4hTtGc8n21O5YArWalbg0C48DjuKa
S54aowTh5oCQ326HX4xQHTmq+YXYcwxqD2reEKkYvCwI3m9fzMgHE83L+XGW
lubLBnR6jOrSuPcX9BgikUShAXWcqw1x3xdoQeNacKkr0FFZVqT0l/8Hz0/C
0Me8QknvjdibPFROakV6eIinpamQ7cmA4dFpZ2HeMWO9DjrNZPOqxaure8cH
6O8Wnv1oIG8ijcsjqoV6G5I1/2sAiC26RrNsTDETwNNH1JmywWagfUqlDCcC
ZqQsuyWOI15SoyujWsHF784sAaF21VxbKAVjiesD7SAAkeYbE1lbpENT3LzG
n4oB7nY7qtflgrm5z/27bOBTyjqwhEOd8n2+mamJzzVdun4uX5/gidjr9WF4
VnWoUK0WcHCP5oiebngPm7aBDFA/gDM8y4WndXXtpPqreRdtSTp0eb+Cwpg/
NHpKqEWPG0CC5KxNKUjSsAMvoicXSRJTlX+zLGdeTGu4PCnjjaEPmD9jZ4ad
HgnZ6UFd4E/bCBEWjbqmdRg1f2qiXsE2PtXSEd+KiZzyophkQgwJj28x6c0G
GsMHMugqyxPyFrmyb/JkidQbn7HhktwfAGXl+V9fj5DbYJlyQVf6VYlaWrpD
klogH4TBB2akPiqT2cqLJrHX3VJhMyiIegmv4jqmf2zdf3NuX+gApeHp+9EY
CXL1s4PlBU05DqWrsiTrtkozggxjj7KBYI41rqQqMCsJ2hGTulJSzhfqMkr6
hTqjusQ7GZljbhlSkzcdw2C+BjCGnGbMjDPVIZyt5ZKpfbVPYHtq9nLYK350
SUCG57K4XIFltn3ZFt+52j5hTboZ2onFdMwhDI5oJkaJvkTvbLCC+WDmqor1
HV8ubuBJ3x0U+jqlAHruvIdR+DFj73xQKAQah0nl1hUQ1enZhV+t4mxt7LMT
GLc7pJCfBsHYOnCMglt8KycDyocewucRb+bMbvFUnayc9DKbFY6CrUTSOzAQ
WzMG3hKU18XNE9QuDiJDNYX4wV+Okda23ZsuvXWvEx3IY24FyA3I4FJd8eP5
OiUSfhnn2cmmJIczJHGWDyLRs720MrkCoeVGWgWNYK2jqfAnRIvImZjnAB1M
gXETStrlPGYuOYQaJ4T6y68IctoPTmjGFsAsSxiyEmLL/ZctBFMzWJlZpIJQ
HaxKL+HXCjbb5IGN/6VxbkBqhbAuGpGcAd/29FG8nzyXJDhYsQXONHYfztar
DTDE/SagxEkn2EZVc4VySBkAHsh799pHmYvInu8cST8ZxapXC5v3OqWyMAne
VotIrsKAN4xPgEJk6FRCpQUd2DXtZbGcQ95V1ifv9jQh2MOm21Pi71nDzxRH
T751dFMw9uUgEHcX8YqIOpoWOS3v53gSRHT4IQfhak/s/iwyuygnc6DM4O4v
oa1Y8VOBuVKH9aCPhm2MUeFJPgML9axbL6wzoQsXMSvcqx/P11CKvlKDjukU
EJ7qb0HuRNZvo3Zgqw5NlQzvdHm8XueEcGd76X8KIHnomtkciANNCtKgy+Jd
8TjdCUURs12VO7ND8XKVP8+5+feeOCHoc+ZD3pMAzGSNGFUM4IEv9lQubERn
jBesgdB7i8T1qX8V2Kt7SgnSZkpr+E5uUiok2CD66+Dor4/1IrvVxrA3V1wv
vHqvXxiZjuvHHASrFg1/PYR/l9p9F2ZIBQ1F26X22FkyEO9lUFgwq9ntlG5M
kvPLqWi2Jz4k/x2zGyTJaw00zOx8vfZFuZrau3E5SqE63k3t6sBEkq1Ju87n
hd8lDlkbb+Ur9Wzw8ZQ3ziIXj9V6/ut0PL0hbEV1q4ZzvigcxfVjnY1IRjPX
ZW0a06qrG4PXcHlJBImttvfJP0a0AMU1BRQI/ys/wFoEIWEU7VZcuDmb1zfi
FE40tVXE6ubqej2zugMJknvfPTn7M07rr+yu+qzIfp+q+ee4kouQzoBHgpU4
znj6Jtx/CxsTlJhmie+tGj+s/JHeriXv0g5kEU3gs4CcrSJLm17fflrFOKTi
dfn2jxWez2mHdKTAW3uQGy1EKvCpWlXwCh9FZjGD9ZyMK6+4VPRUdhOrxQ3h
6e+Ip1JVoy5ZO0L9Xw8rONJA6//DO/UUEa0GhmZSehgjSKpDTvxNRUxthiCl
waGUkTKATbL+d0a2ueGr7VqhoSA4EKJ6E3PMxP1kIEdv6S0F1RrJXg7JcAsN
idEqrY3J38eTQCd7RkvW1NggnVQyz06VUH8h6i9YIWzNqDJ9A1zxcsVoxDSl
KBzWrZvJ9Cj0ep3m4Vc84mxtrjJE+Aeter38NHxMEiDjvAKmpqOWO9Gp0SgQ
erVbopCzLW0=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "OJXsOzX3SCOyhcBXS9yryN9cWQxQkhDHUr4mzQikLKNKnB6JkSYY9xNnmYkvVOJ5f3SnsxLM71tWjwpqmyTCVkTt4jikDmXDCnl6lQn2TVy78ivgbebFE/F7GUr3Z8AASPmtz4v12cD/Cz7nTJMTG81IGzEoV1S4KsV3MBcbB+1TqTshtjzQ4oMMPpNw9ltjOjjqx8CktvtqLiQWjnKfQh8i3R/5yQlzObBDq+VCqANtp3J7yp5y22+Gqzr2XdxPhhqdWI8am3cUX/Dd61VOxRjTLOoo/W3bcjWpJkKZwNWbR8NnoHZTDEUIaaMUZngVX793bxMVF/DlIFYHkEXgfiAeuJaPRuz17vw68dvasrwdN3yg8btkqN8XZ1XMbyGxNPPBR93gxIpzF/yBuEw9Fk0Sg79oFJ/QK/Ju08ES30gd3sX9p+6DiY0U70otzVbtsxz7scd0mFmNYMYlWs0LKKfPDKKOaqoSFi6qoftsh+49JcWn3HaMKOERzBWpeW8PzwYnGWtqJLNSVVvEPo8IuILOL8fEcwCGGWteF5Yc+qfwYQbbqsqwXcqDyT8DH9q2BydvKoLPmLdtopwMaWbpXEh6b9OCJq1o4l/Epqp3eaR1OfIsygKKDRCUWaSLqnFyUKre6SZvgyb55RYfdrkrhpoeJSEHNNinGPc+fClECLDSBsGRXGELbEC2gSExKZFsdz9u9OenTUYJ4fye877qjoraq8pDDCuq6+GCzWVK0ue5VqE0huFI0K+yFXBHXQnuYIJ2A2uq+q50G2kdbqVwP0OWxyBlbPvGtYy/VhuOhN9O4pilZl++nZn72hmDKO5H26+Dh3rFYPY7SlrU5drXKwxjeuyDM/z/964/Ws5A4N3xLzGalFv90Yq7qEzg1mEoFXUk83Y/8S6AZSZVjaGlxSZiEiHlaEIU1C3K0O5o2N7dDVyvWTzU3dsFfOo9A8ND+CU8+UWpvycgpEkDQYBkDnp/AZ2qiDzZpOj4upBRHlx1to41kcwtQKJluCKaO6Mh"
`endif