// (C) 2001-2023 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h/OHrq9BJgoBIugx9YTP0El02dGgMWBZB/M9OJs63hBzMfThHN56XfhmoIkh
OQrxMaWBua466B9BI7x8wBacZXwoLafLhNYt7ufvlc6T+IcxDWQGHiQZMfS9
44JuyEb4HkJOXfEsLLKLkVUuFnCOshb0oemnkqca0cnbmsXSzGdGKGz8heL9
gj6FZeGTm/L7uAA40mYC7zpR7p6WuEnC7jvSdjphPcXt9gzVQHOoBzBV5CZf
fEsZngm+kZk4nrikhm/iXgd5mp2DNu1Wi7JBkJmpAuO3I7EfGHhVgYlWo/up
nVRTIM6p6VWKAIo1FGEm9TlLl6QSobs7BgVE58AUow==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jWTjK4LYj9jBBYkc0XPdWMwmXiIbPoZMtrMtBmuWHP1Xk8rwNJc0ebDWHSJ0
ibmo7PfBSV/15m7f7O2lG1TdbgbsFFRvYep1JPwsqAQSmhBAd/IoebeEvIp4
lOf7PV2r12/qD8bRPML0wqacZWw2etsRfRaxwAnGDYi6ElfIEoYdCf7NKy3R
YQBHt+wHo3xfZ+yO/GA6MQ9SMqlONfiRz40FDKZ3MXkiPzXcMjvWDOienHz+
Vd1RWna7mK190l3jnEp2vKFLHuvAsBL6uu60pmgumRymrdIr6s7kpZcN+Ft6
HW46QX4bFK0b83tg9SQMJ2xBbuOXKC+VtYLtQLvCkg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Q/DHWm63TrO7CWVN6WJ2+nWmvis0ETVeBzqpJBpWoMfr+l/GjMiBXKiWQ4ct
ULHBNVu8s6wdhuL0d6mcJYVm9dGMqQdu/44M8SSAwDtOJwC4/4IuM63si41k
yb0/Zrqf9PzJEG+BFz1j9dFifYSzcu+/I1vTVLEqdXS8n3LH8ukky4mDzniu
UDIyUzmoZkbnGP5/CtchZf2BHfsRLEVoyCDoOsbkah2dnd/XRGqEGieYSonk
j98FJYFurG7m/Xd+wir7ugFL5f5oI/AP2QNATu1ouv5SyFQMEVEw80cvfgtZ
S3YoQFLB1X7gprYoKB2ECk919IBudhiOSIvV6SHYhQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DX2o6QaTuEW1ZLsdxXYDI8gduKlBWxwiMXjLG8ToZnwCwrkjedVw06e1dpO5
0SSiKdMhbrnqs6YlxDPiAiEN+f/eImlVnizNYPwJ54lbU3mMaoqXEEflRqEd
Wi/+uOPc0FXodmWDGCnqb79Gdje45OkUUcgJI4gkT4DeV5ow13w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HegmvhzH8jIpQg1Jw7H8aZpMVeUr3jX9rWToDKRmAUZaBQhKuACgCpNBwbGR
L12Ub2qxwVuwF/GKY9LzhYpgmmrZeCi9CTpvK3mDKpvYRvswHUIpovYaprkG
LOQ/g//JnQMtQqdU8yHHtlElySMZynhvYfgKkEC+m0CmAx+CPsl1IX2YE29w
uKa8fjFiOh3w3FXY9lO270alB0ZwapzhemnRvBeeFXh3IvGQnmgmXgZX/G/e
pIljrrktpWBsrsCqkPOMxenxRn/DwD0SfsZnq2R3sFFgNz9a9fV68KNaHdqn
QJmK6o/Im/rwF78pZVlXDUJo1QsvGvTsWkQAy0PacVRhZkdRx6Yza3lg6phI
a8RBzcI9WNi9bOGHiH4Ten2BePwmVYYSceiNRyUs5lhpG3FVVlYZegXINypg
/t72mnQGFsWEfbEOjj2Sglbkzj2/xCmczlRP6p4K2tnYjxMg0qjN65aUGYAt
O9pWjRjyzWjX/hfT3eMFPQcccWrm+mVC


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ogsoQl5FkJnsYzr4C6jcViYEypBqketyXZDygMqSibAmSJ84YrfmR7xdTybY
vCGu/HhkqWi3nzQkkmPr2DjXigs/D0zZ2hGEfLsp8USeK8go0MSoNCyXh/ji
8Rxh8AdHzMwxKi/PfycviQQVvfG6aSaUixKLF/mJq8bIqCeW4Rs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NWdqnbJbIk5023nVsgR8fvyERipK3Vjin3A42E9u0jq5m4ew7E1PFwe6UivT
p22u25/anR25Imn+OfiKDWQiMiOkzfKrcQTYH/Mww8FVbgW4122wn05eUvoU
zsuCnyR/qCeOfmfozYec4HsGBLCkYaQ9g8hmIptCXeWjMjG800w=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 38960)
`pragma protect data_block
iW8Y/seaStYRLrNNqvZyiay4TLKzPZfX5Jj2jciq38x+sTz2f2W//2RpAdu0
ESEfDaMuV5hYgzZdqE5R4648N6qqva9s8AKX1OYb2/c1cDloVh2bdm05sOI9
4ANeXxM2imrdNkq4f/q2BPDPQNLyWVqmoG+32I5hzjhC5/1rRVW/YyvHraQF
M/7wt72ZmrhVzRFPMB13bFmje+RbTTbPQy4dY6LRQVDZUekglCdcwLvhzNOu
ah+i+IVh8C/16WSOKECIaavaDSe19RzZTsjOZc7gN3wlcjK2XjmceVBH4yhb
OSQgScQLGhEBsToWl9fUtVXMTm4ydztgLz26i0Ew+AR6ug3W4FtdEaQHkh/F
9cdaMHTUFR8ywxDEUJtvUorx/aKrN/OvzH+2pu04PoJDiD6BtV5LUmnjIslz
pye/QYHtko5uNLACzccob3By/fsrHJlk4WIi17uz+PxMiH6UPmP8vOBKIM6F
DHR8yG8bSd3yaO34D1LPqVAVMKXPR3J83PPfM8wDEzgZptkUQl82AEZ5MdVV
yuf6vMhylRk8dj7pIkf6czpfzvLb5eUJThXA9lzxvRJJoA11BeEjTQBQ0uZu
WfXoImOU6bCpLG2M3LK6uvj4YCwNBjUWPf+ii0KrnOaZqp1nz7R+sVOQnwfZ
+ZwsCI2VJAE2P+6Rc07b+8EqFisdStZ4IY8jfj0Q4RCjQfCx+xky56oYVAp0
gVGqUlKcHQafgMmngoCpHdWmK+acR87VjTQYm88AO2//HDwPH+ff//TW4/cv
7WD18MH0+qBu95O45+md3AIbKDtc9olNAA4oTaqtKIfbLfzvvfMXBy/P3K1H
H7FNtrIwOyyq82UExFKma8hnGEz144fjgQgSVZzS8QotMGef32ubUMGON8WR
ONES2lmBOVA6PBWmmpGBzTfOXMEwHegtjNHGqm/Cj6+Yezb0TuMnjfQhasTJ
1/4W0LsjTfnUC3Uwcd5Aemkf3GrsAxLL4oAbTG/8W/3i3vMNX3REGsX7VDaI
ME2EuW8jAxkdWp+0U2D4MNMgH7kJcg6RFDrLemDSUyOTh4yXaMcKGlv0lXeX
GzQRC0L9THYWBn7NEVI9I7KUyHbefOTjW5rKgZf7e9rvi6Qp0dzDC9htzNQI
5s21S5zg27/4eAze22XjLrIjm3ja5l3JUxsyj0l79GTTzXwdSR7QKofuOV7Q
zPwojndYdmK7pvYbF6yi49FEnhTuA1MBkOjt4My3Brn38Z6i8QFC0b1vgAVr
XzmG00EAoB/d+BbfUnGkiOfhIuV2PWNffcYAFmRm3rrHLd8+P0IAhsq36TAs
wP4FsG66o1v1W18OaGgqDPqOvQNYKLGlV4GGevdMEX2+clYX8+lwXAaUwpew
bW0ezOM2Vp/tn4cte4B59oeW7ugBrN3dy2EmCG1lAdZc8SIgbXPutlqwfW2z
EXjd4fOwpWWIhEdI19cscev8784hN6CzSrYJ+2qXGEioSAKdmQ3ezQAABxpN
LsRr/lE/2vOQh7HjqVzlcGCVyBnqsyzDNuWi1DC/2dk8oqYOFbjmZET2PmW2
blXdOcbxRUy4cOEzG5So1myDXpkRp511/wG7uESAXD2Ggu2FgN3hYO9PReZC
O7kzs2wiwTQZPB10Vp7jk/bVZjqXhRfinsYzP1V0Iu67XNLbHvycDXjxRHHy
Dq0mAFbgYhEfsnGv8YT071NfPmPSeI1wnhyl4q2FPIaiYJjckr579YVhrlOk
60DZdr1J1eP36MwcKErss58iN2w7KLx9W1/iSmSFRG5zcQowVru5L+0C+nZ8
TsLKUluoFNvb/2nUBgLiERonaPzOYNNAUYfifKpLePuAMmP2MqYu38VxebOf
XoesaXj11UgUAG5H5dX1LBsP2ZwM+44LBiG2VJKw0ULqm4dhLVmNxH1Ifs0X
rksnyfMtWpU5t2wxF3THwW7bbSQnRP+cXj0BqBSonN103oEVUv+lt3V/zLZH
NQy7jMRGhEXxOih4PRabcB4y7fwT1/6p9GNm7lPk3l5gFLMHSGzZiDq3yYWL
zNRBvKZ6DEx2CTQLSvKJgyIzOescgT1cGBLYT40UyGbgzcYvTWVIwx0q3+uW
fMQHE/PVXvEYA5JI+BslyjLQ7Vf5fcGkM2/gTpGbH8IEjoYrlc4HrodmPeAV
eZGAktC8JNc5p76MRtsYKr6Qnb98LTRlaHNIW8uapZhMvIWDvBO6kaiEfA9c
YVajWBZ/xx9J0J80KNiKIDeQ1ydDEQFRfKTD8ZE+Y1b7z/dPJM9DmKx5v0Yl
xqp/g8sgOhgZwautKJR2fLZg8FP50VshOUMGlxL05zAOUZbVahu8z0FDqFNT
PoqNdqQtKwUDMDe2zwQK43bC6tQBLOcYoVx9GgOaznBrhdjnKDeQbR9XWLXC
vY84jvwthYSWYP6OPfOSznbyPJ+vamx8JqHeOPRARKMi/HFcwrlgCal6twNz
ZNisKWvBsk7G+u3WqML/SPaWFiAFd2l8y2cgYujUVpXb1Oxv/Z+yEZD1zjPH
973lwe0bk32N4Goh4EZFszS+srIgZ2voJP/Q/sB/qKEMDxky5kG1Cnw1wJNR
VJiud6C4yyLPaSG4j1emTFz+9ns2HMKa4rQ0J3rTAeDQIfHCqqV4nucHjVeo
UUBlbvPlo8ZD39l8GYY+V7cC6oorE8W+0e2ivEEPMkc2oGDbDPxP9MLdwyhf
dnruQwjEdLqKq0TmNysck1Qm+Vgx7060c/DjHW+//4h8b4mymCCSb4kCi2KZ
eKY98KyC8VeRJc83poD7YiOSs74O6VEFvff0DToHu6JtWhWNiE0CnNlKSi3L
Ut6Xbqay/oQ5IYCENnTp4UIJKVN3HlDt/jI6xwW6XtMXoMCpUpI3XBb/ziW2
RtuxPUjy9y7IDhewVVD7JmV25GV51vENLIMDkoc2F1irXEIBCp/ayiiqw7Kn
Iiie2ddPEZRJgg4+Bev3Gfn/7Qv2z72LYouDrG0uep0OY62JA6sQvnoB1pCr
g2bhdWYVT5EdJmsm/kpo1YcloHkjwkVHx55Z/47OLNEi+JjJinvLvH2n7HHV
STMkEm/P2T3DUSvp+3Ago8Q3NR22u/ODNfurdNzZ28GbwiaFO4Ja6eCeZUq9
lRaBK1ycSMLR6wCuQzo9HtTDHuuRB6Ec35/WkUU8Vg22OCoMDR+P1qdxw4wW
QUg52nustBVlr0vz57UwK26lQpxB6MnvAb8GqqTW+qn2JSQcTmMLb4g7M/tM
HRoan/XtF2bEctaa04XcLTNWK+hbe35ZcrbZUQCgcKgKttHK45hhECq4nq7o
KwbJ7KAJvgP+HEDJO8D2LKOqzL+AK8EUFzvFSB411foizdidC1lBhiPOusBF
CbM0L93Dywq5U6uqfIdJo/l+5ENOLEiiNwL3cLIZnEMU6ZuRUJa/nM35vTOp
uouSLfexv16HaUiweo762pOZwsso0G6G2bSIe16WGhUaz11syDqGXY9WEm8j
1Go5p4HgTKkZYMTTYFrYKPcvl6EUDrNSqSJ+hDBB3fus2rpb6qfPDziSUwKX
KhLmKlvaM+9ozgjwKQKTkK3rbiI3KYLVZ5Y0oWjOw8/3FFbrmQ0jX1Yr69l2
jZkPAL8soE4U5+KXjGrZjFr89owocpNQ65L7un6GwB8hzCgCXQ5O/JMzDns9
gG1/ZobbQyalvTNECCYz9yInk846mVZfysE8lwpbZMVToQf7nnwwR4Hjmp4L
2khVYs+hdtJbOWs77oGre0z94SjHFJaeo/mkudIO2aX5YfPN5TEQjfDIDjdD
0g2+v9TlPopLCkHpX55IBE3eTOiaDch0oWrye3hOhQVjGD2T/w7pHhg21Hwl
Sd2ltqKB33ah6iZmsr61kmwewv8PQgkhJy+z6z2zz2J0BPDO+MnM3hhnJY0+
Bimp2as0yPgFqedWIq74jtq1xe6/iQisJGPwbJSU2MdY8ek02r+JnIlniZqI
HELdFNidWvaKZwFl3fhbUpD1nBTgAM+/s4SnBi8mEROvK6+sQoVddXrR+hXA
W9hGwSpdRPYa7zLCaYQ2TB17rLP09Ulwo76b6SLNz/pCJeQhdu+G7OVy1wXg
MK0pR2NcG8Fl8uLbav61TJ6m/VM2ipCGbEAbncpw1W5JJ/4ZyhPU5s6J8UZe
gMZABL5E0F/GSLngqV1eelSvgLdZoTpnhbYBFXX/+j95bJ4YYTJV29soqt6/
1x3hhq6j24d5GEjjL9ebmKmcr8M0WQpZseJhSpwRUeTf+qgaTenYv0RytVFB
gA9I5VhdtfZQgnUZvnsmx3XCIyVmNd1RLZGHHXdjiFFx6beSsL4qJzD4+J9n
YnORJOt36nOYONpS1lMc0sVxZlv0S2q/rGwiK/r7zPpza8hhpiz9zmUYCYSS
JqBnkFfrrJqtfiARFCzJNmCAYBH5kVcn59nP7/0Lzk0/Rv3ql2vkWHeygT08
q0s8US8VanIS4iye9pqO30BiCyh/JrQ+9j9WipbNWaHTPwRro8YwqQGGpWsi
ILx4a9R8xv7/hh1tXZTpur1zockgFyzgD5WEUm8U0NkyG3n46f7rvyzbJyCe
q0pZ2DweQGMuW9t4hnADbeVAREWuplL9zBNTzWmvcbS158ez/pkSTGTaFIC0
HDjb6Ao7ECg+mLHaP7kSoRpGNSnV4av8QmoYwcRJOmTxQaHSzTUSYlX8DfFx
iMzUvz4hyrEjs5NXeh9RSuPgDtk0GIK4kmnnx9xu2RhHo+pw94WAVpC8hOxy
2m90mSQnFRfYWIPJKmQUwdj567E3yqCXgnP96UX7Nz0HOpdOM1m4ONfVqPzr
2qbG8wD5mvX5XFXAgh2QxnC+MoAp5/vLtR6rpbYBxKlvo4wDfQgj22Brbbbd
SOborYWsVNoQ3YK1cdLsx4ES4o/ZIjyq/924qeko6INpSSU1vGz6PaJegOhZ
LvTQ2KL0loxBJ831B8c7LdD8iZkAyl+xXBL8zjb1LmVHn8+vL3btgp599tUX
M7basTUuWNLOOtBhZ9k5xl7m+p6DfkcpGanHMZYVgsGrnHd9ZHx0/iXfIBW4
U91aib5ZrVBOwBuGd/1AP5eqh8VLrTGmqGE1ijInYmTVMBlNhV4aUknJ50pZ
QemKTZMSxATXTfdkwLEfVNRG4PYzrK38NVRnjEUFJAzuWFeko0nDokeAzMYv
JP4rE891jGyR966h9hAi389wNvIjzN6RDQ1yZ+aYVuUj0q6eIxSclnt2/qYZ
hlDEgUMKRuXXMObdLhynZpPXL5q992fgN3l4h+LnAh1GuTr4nUecBC0Q+kRK
ksaTm9RewZtdTvTxbx3EOgDHIC+aWhXYQVftbGY77h6GBUSgKCa6M1jB86I6
kKwqjshVFEAmE9i2XE328qDb4IvM+rXkN7Zqj23d15p1bpVsNRrEO78M1y+j
saUdirkSrQY7V04ojbPKucrnQjDSSvzN1lwzXq2jORt7mZdjZ0ISEgQT91tt
X9seWDw70SR6clAHkJh7Cdgg20AvKI1Mw6W6qDRI+7yCg8V5WJgrstp07Qvr
21ZnFAKETLXv/hSt3JnWg0aZbC4xLXnZ1dCC5lhio2oAKtrcbmQeNHpg7vWg
iLaTIgKcFK9quod5xMwRlsa4sDLXC6wlMAd8HsEQ3nV4eyw1UePYXzXLfGO3
SarrUudY9kwgUjFAi7WKlFYJAZbb0JtXY7dhCOXgAFPcvPXjOvfNuxPnKtJI
t8wqnqC0fuWa4rvEVRbWrcV4m1PixQA62rAtxMZkQcOhk5zlzj/xMd/k39Do
A+WkrGdfmdycGsr2Ecly1DkZXtejgmX5cTgMzgZfGot0suYZXAa53cZHXYYG
jnx+0N8r9ZepHI07LRnm4/S5wwYpOabq8zP4bVgOxBOjFViyd6Hen+JFpEtY
2Tm2vQ4OGJDE7ZllBeRXWT1XYxL535Qz+okzodRUljrf/20i94mry8sM7o/2
8Csr5mL7V0FXXgV5O3+Qm0UXRhSx+YTozBqLc0goc22RX7APsrLJYWNYRQie
OGVKnRdGVkPBMGChmgIZbjB2cnE8BvCwi3gj9InmIyx0yYQUpf5BudrY6i5F
KIyqohAgCIPnM1y+u/dP9zaNXk9Y1H9l8ghgtO6tBmlZQ6bUXqKwY1JBwTSZ
YMXmSSqXwUok3OT7O1n0Q2CZsrN4SOJiWypelN+PJyjSj1K9mL9sMtzaM8sq
IszirGyF0D6HQ+Qf6c8VjPfPbd/Y187xhDbBCmgf1KVpCR2QTJxz1n0qYHDb
St4yzp3S1bCEmQnLD9ktD6p4X/sRo9g5kYuay/BvM9SAQMQTMIInWK5Ch0k3
HljLM23r6LwEbdZBcSXNr8o+UuTlo+wvCnTzqcRfsa/kfMXn3qmiNQ212o+I
SDpTvFrwdSd0Zp1lVtE6HYmmRP29BksFhVVhGJX1Kdzvmuu9rIMUD+5V+dMP
kBMBXu8D4zlyBKK0Jbou5mdTNlytrbRU2fHEKYvLDKyzV13iZELUPX8vixy+
GCsIc8Vf4gDG+J2ux8G9OxwHLFxV8bOugOA7jzyMEpCZlL0CPjM/AmdhAr41
cQe6M2h0xM20WmJIeG8ziV9bWamhRqpZtkpuJDhs+js6ifz99fDA5MPwTD8s
s1xhMOTBYAHGL0pu5wkeWoJP7FMUxGHm7iGIf4OKRJHmVumGQ5HthD2n+dS8
Ci/CK5YxzrLU5WE05ZQExT7j7r8OnULdYnS42K23sAnjEm4FGD7taEo3FGo9
QEPoWXYpjQlgZjVZqQ6yVJtR/2cUNQ4FCdZmtxRZ15DeDyXAvf2BPyQRfyJn
SjcTXxO3Td9vwT26OEWcfVDH33dLf0hky8ZDnuXxWCdDwjZbmKi8QNJWNiO/
hTpW0k+n4tJVDy5WDiZ9k9wP9f9ZMhIPLIB3+AVbRaQcvcLVwXfd98sQ19yb
zYUu9n7vuRERt2ZWpNg+wNbeZcPbG12C1HFjDR5L5Qpt2IH/JTNjjJ+Uh752
qc7fF0z18M4oLMnr+ghNzyiCxNzTa9JsnK3K7QkwMN2y3dmVeEmM2F12o49j
olO4NfHb7eRDLFA5IAGg9ay+18AAwWNfMD7EfAy8QXnFDFVpK+eeN6kH3QBD
gn3gl2HOIB3+pZtMD+qIptuZ26CkEHVhfCXxN4gisRnI+YSHUT3Gxa4Mh224
CxEvtbEnI5uivR1Kw4sVGkEtaWrJAngeECWqIkzKg2P1WSxJKajDaBT5pI/5
jeWREUKfuD7djY3BamZPDXwMJwrFZ7eeV/EfaPTDGiXxDB0TtBiHi9hLBwfG
M/DJgzKh/nzKJCsssIlCMdDkTzmqYuiX6oFQeM3xRF8Lt0vawopj9PBSXv1H
1sw+JB3fwyGLkh/BSUaBLNxDA+YLTI1o/X/LzJR2GgCMuPy8FryeON9isfqS
j2WqxF5JRoUMww5yMdqQ0A2AQEvvDZFb638jNhsgAvXaqOpsNl9g+KOXpAnp
AmGrOfe+lyS+ht+3zyp4Xog3M0wm298+vw6jz0eAw6BWYIO258Yi9LRHmbZm
zOGLgxtnZ900VZISaN51yh1ttzQMOXSTHVWvHf4jdepKFZHfsIyOuntD3wJj
jJfVDcyoDmN5F6xduWcB8xwjslAELCwMFTJDXZg+tONSrLuqtSeYyxbQ8y1B
RjGqPqPmbg9j2ZWnL7OFFc5Vu7uJYjxp/+JzAm115gvD10VQtRel5RYBE8xj
RzWSqZhErXzP91o7+fN6Z7IgesfWUAvqgXlgzj/Jy+YST5hAzrG6uEb48Xpm
hY/iMY+rzhG/Qj6XnA059IhywUhX4k/8vtVOU1/3l17Y3cRHecDLdynoPExm
UMH2JMU1inH3v6y6KUBSw427ENiaTc60rn1vbJhcTtF7Rrjcnub12Y0Zvi07
+etQ0X9aZbFF96ULoHyyftR5RFwwdEm+JWrMC/PBJdNnIKotBYpCyl2M/O+/
XwloOd977Ocofk+B43bTFSQxSPzreNa7PW+pSz0Jpk08k4FSA+GSY+Zlma3F
gEVNYlDGGNmZV5L71iH14440Kt/YcyNrS60HdIcT1gHrD5eD5dNQyitWj4di
UeDc2kBj8WeOvTbP1+w1uHT/BKGA0prC1FreuCgRvsdZRWnctzlULPOv29s/
Q/mpOIb3tmAc3KFU5ZjECZtVF8Raww2dEZFmak1tOJk99ic1b0UEzy46mMzG
XFIuEcdVARjzFwrceu2Iripd02l5F5CufEH8hW3EGDyFQFIE1QlaEEWsOUD+
Lm9V3E6fa9j7h//JmJoxYC7biWTGmdh4deKkuN+UTc9E73DYTGa0QpTKwnU1
d+tI6vCU7/RDT+DTW+TYnPbXnxZ7eia4LRfmFLX9gyG6DwkSQWeqmYDxswpW
QFUWvRHRoaevoaEXePXzJ8IyzoDPEugbhaGuAGkXi6Nud0Us7s+UgNnnkFyQ
a0RIWBXtedgZaLTaUb/q692Q+0n1lbAT/imlKtSIpaD+jNdI89yN3Evp1bGa
rUYt/L83AGgGcs7kDS1w6xrVF2WD3f13/h/rGP49ufQtxuU5AVGj0clxVM/f
aUPPCHaZPihoFOg5AR/kyV0kvx1AG/7DUNWnpAXRD3+AzCnd+0Oe+3zXwwrM
7Xy42pg3NdvPYsf+QbKyQf52oKxEPc5VQP+hIJkhT4TPN37FJRZS2Gfh3ceU
E1r8Ca9Xi1cYfsQ4iRWedjhccUMpt3QTm7lfSKwpJhb1ZQqNxz+TWj/GXhRx
YV4TM/XHBG7v5GdBFR550GvGGBYjmdiyKFM3fPpjV3WJ4yBgBtIkJ30J9nHu
ePMw/Hjh0WhLZXnklHG0uREu/V0rFrZ8Z7240wAt73MUCTug6/hDM59DR896
8cjElaBdSLwO94l42rjwpN/A7HfBSZ5qLAl9pPS4gHpGOL8d+81wqrpL9W51
18BNsRWx9h3RKxyTLj6hwxpffUebw0FX0qTTsrXl+QHg1hKZgTTE21JLRY/D
SQg++ldl+Q/F+9q4ybXEokQakDmp8fPK9H4fIV6YCiyIqH2nevE8pLJI1tzC
dQnf+HQZWrc/lwhsuI31lwnvvAt0HJfF3EDHB8rLLkwJFDaqTH2gTqIvs6Vw
BAMWeXjmcqn6rkInhhzWufKUr240lAWqJRSI/+FmCQOvPW9fLmz1xYp2aALr
imcjf9TMiSUuM4g9D5HvylSLtYUdGiFy5Ktjb4ABxQxnz5JEqhOwGYf/18Nz
xIH8f7K1XT8woVxb6CnLOJypJNJ3fAxQa0kmx1O9hJaji8tytllk25isLwwd
i4rlBTWOiDEpxjS8WKGJHR9anlQB/hFsEKh4ED1F/wNdGDEVo5zP0cheXIs+
6AEbipJQRRi8xmCNQKbMLWOLc7lKw35zl8z8xoOHVEfDQvHK0ik3xHNbCxrh
yyciS4Y46w3vl0LNOIrLRC9KzfgTZNm24KUt5DTj6OH5z4YOWoj9OVFg3E5+
/WCgnIF5ogKufNO1NdHJj65MxEmxVhJndPbNQu9y1BgfIN4cO4fZDdJOCDvX
i+myI6JHcGvyZWJ8Ce70FWnUB9TPwL0TOTpei4STzlmhMnVsVd7v8t3/bYvP
CopYbK+ewKULL4X2j2zBsKKCF3DLvmz+/wszMmdMOJ+4fOr3Jp2Y2yIGIaiu
2Izv8yES0VDkeuFoQD//0XaqOnuzVZHLOpPq3mmx8sqz8bl1SjGKyBZWzNV4
6V5s/O7V+xzWeJjMSTmjKz32zV9EAz9Sl9Sd+Lh+XdiRev3rRQatj59u/2eY
z3tOa1J8F2sVv5h4om1HrPnmoNsvOTSB3cKjSEJ5KlrG6KmmT3KHu0IH+P5b
nbf2uLYCN/lfCF8Qr9iYwQ0a6mz8PqEGkFZ3V8QpB5Yt3cBVi6Mb+eiIeI0o
Zj6aNn5etU8OPOP9/bPpqeTBrC5hLejRQPjpMBFHzzn0hwKNwu0xUId/n++n
B7vMaIY/lk+ldAjE9wVtYc+DR1otIrOWxGGYVID90WoUCeTWmyvwpQgb46TZ
d6SXTRMlCMYAw4UNYcwhOcMp+1imGTNfOYnVTvd1A3X1a/yUZNd8EuDHSTFy
nioQHsJP333rWD79Wi+RLVoksypIbOPdb7MCAU2D989PQllpdDhsJ0i662bW
y2TgzkGrvz/oySoYB/lrMthnLgIV5SRDpQdKDvWEdeJTmJRkMcv2Py1VJM87
2SUGbcmPh/HBmRMJoO0JaB0CIpMj40tPVutrJ/TLmnmaAdMOFJVHAeOR4oVb
kdWt0k0NiE9vaa6kifZK3XD6W+/lSBGoYv/VC4NcP5QBziOXh1GMeER2Q0c6
y0sbUzHBABFtKasLYpVSJJIaBW8lSEyC0pW6VWm7t/HheW5VMpKSBG64MPg/
piQrnWM70zRSsNT6JjAUEa0DC1lNOFOv+PKcQZ08tVF9YfJNlts4GfCo3euQ
a818zXLdJZengMyvnaZhiSw3k3aR6ZSjLEvJlpll1NJGah+Z6zGiJRPUifi5
qSyJWvDGREmb3zwWmyLxjT44TR1bERLCxZ/fTTWYbBmrHTi88EecVhZAMbrU
fw4LNWObJR+EWuYMzHZXFa58qCLAIA5g6PHR1hzpUUdZu9rhSknTL+wLG7hv
k/Nbc4z00y4GOoqcuaz2XrfVURvnAaCbE2PFaOaDGbeAUC7/zJO969GBE/Up
ZCe4tCSmP5XnEdY4nRyJQjbpC1+fb6PBnJVbA5kiw2yiWsMSZWzY4+VEpJE6
X7DDXsXtXLZGOs0d05NhLoPwYkLR740sH9q+FKNlZ3w1M50KmilKd+EgqGN0
YZx5uy8KfU1Zc7uM5zDEvpzGDEAB01H2YwgeMHZOwG0pPFgDOBUkwnrEAyd+
7NfZxmceAayeaa1YJuu9MylFCxdzWNrzJw8kzb5aEBYTtpoUYqgNEis+IqDe
Dv/mo59J3LNz4Clxtqgg4sq10UQtNnPuJOkr2HwPlGLpEuRhrlApRgZ3jSQc
g3b8sVcheLmkmTQXQm7rQVOrlP2/VNOTGISpCunTzWlS8rt43jm1KLmmP0L5
xAFQST6OYOTZ96edAiMWswjy10YPKZC+EzqpnoQMqH9cT/Jf3AKPFnza/vYP
AfJsm7F4prsMX3nwO77V7aKkAiQkJo4ZoZ4vn5kDDnPpopv2nBgkspRvMqyU
HNgnoqx70LnEP8Y684xlYe+PVz4GEl9+IHTZ0/Efv4v1QMVd1LxH8z9/Dr7F
hOy/v4cNfOdQ3/pQTHuITsokRzTSbIATLv15NvHCewbnVHZyLOoyiyeD8Fr6
qH2BKk+plkoh8n1n+5+tLYKxTLvqXtKHcGPdzbfKo4fKf0U5/sQcPilQVPZs
iM0Bjb4BoRmQy9I/NL7buz3lhGET4Tq9+m+oLkwbapcLt1+3ZDKh6rJFGgOd
3rcgUtMRDQcm6hjrXbM8q7BphMKScVQvGU5nddAmmaaFYaNlI2MMj13BqBGH
Bf4wQVKmrumlDM9/Oe+hR4XUv/2ajyYeVMmJq1YP2kzWI1QYrmS27N5UWRNV
t2pSXqI/VZB3t1qmnd5iJS8lGlDUxmnjEVtROro4NYxm/cUxkRihjR4Nm1rB
1UpP97/MD4fYCt5ODfQ0T8HRyo7VdRj1FT8noKtxoCRfOMLiyVQJ4U/6lEv6
UJT4Va9i2inzN5jLlhK+fpu1J2DYLHF4fw51hZlvm/O1Mw+BoS7HFwHV5sip
mpYACKEmMbiaTM5pMzGsHpeZlVmxpC0+RxjHjRcQex0wTY0aOEGTDhn8nWAc
7OG4W2wLdr4v/EaGxyGNn1NTJRM4CvdGqdGPv7ueecMpHjUcjcljCw1cLbHV
jmupCsIqts1odz4ViNuYgt5zvLjnwNYxFmL2jjjRnMHCyahmWy9yDWh3Uc70
olKpcOcwFZZMfyp5qLRM6z8kPH9mSQMUjXAKhXTSciXHiRGuwxugwt8jvgKM
Hb1GUzILWk61USoVZrMSrb3GWQbkNd59cI9awgfBpSrou4dwpuDrJmQnPdI+
Gm77uhyyVBCKP3G93BDJaQI+fDiNQGd8rY9f61zoLW59bSXbZ92sxjJcFKyG
uvjuLf4H5ioRvYE5+mwK4ZO7u0DM6nQld1V6hGDknvjE1AcRtjo7LcjA2bP9
HVm/FtPRrwt+c0yydYIkKfqJBzmcceH/38JMy/Kznjdpp42YcwgGQMVL8Hb8
teQyeioBeWs6nVpBjk0cQkI1ZoV4RjDkJkUW3f5LoRzK5dNNFe6VgGYWiY7E
xSSPjIbfsgtbjX54NaTgOYvZtPK6HChhG8rEY/nDAnmq9zYieJrUkms5Pb6j
5JcmaYgQvRDa14XWGsMOAIyfswr3jhp599bWZAyGYrHRf85wfPnhJTnCGSPR
+1x4dv4AYD/1V/IwjGLyWMS/0//frKu9ColgY4CeHcdeFwMauhwNvopxLqVS
tW2qq1n2TsyIkyYrWFdjQuwxlWrCC/2KrI3aVFmwJHfL0epsjaRbsWWUIeGk
P0Ke2EzIqlB8FBfWDvzkUMmwC9uhG5CW+EzG+1Rv/sL5uVk6dOg60wvSXyhG
nlY1xW9Ap8gCV1oOVM6L90jpIbE49ZLMPhsQeM+FBg2ugx2WES44ur4s4NFW
x9ik9CV0I5IYoF8AtXzOijuEgQyEk4+vGJ0zrT3hpktuNBwDrUrb4OWloy0i
s921MnYSUlub1sr61RsIyBggYiH/QJSz6mJt//ITHtnELmAu5yvfjS7grfrK
mG/ERpm9SluORVFeG0V8zi4m+dUumEMp3paIeEX2XLcJW7IXGiN6HLbI2fbF
ppZ9y2TgDYGca2J/VMr++eivdg+9D50RZEZn1PvuzUiW5sHsKk+DlxZUGNoH
/mtAYJ1eMou55F/GNGhmjSUo30eSaJHYUCGPMi8BP6RNGHAivolyryCNbfTp
dfBw0W2reoSubhkJp2xl2WSawg33TS8KBOsNmy8aBwEnm1i6FYPxqbbucnm1
Ym3S/SfnjoqSUdMyf3PwNgZHZCvqVYpnpulbzutmFzsYoVzD1Fwb8CCesIZW
CakYXOQtWVzXg2qLo5BsYtm3Urq4B3FpVHGlkTY2blIuJwZPjJyJnOh////z
01feadYoevPev/Y+GrTvfKnEk7LQZ3/U48+63DowbiHVHS4TYQHX25MabAxS
Ah3v6G871/4lzPjfPNqdhJa8dwJbYcVfSjbTp99Oud5w8UZgfF2idtV768OV
D573fhtZueqM/t6pO6l4FZkBJHzP5S0ecTKztzTOyfvyaicflB2z4KrBvA3o
et1D3+CPKv2nuKrWyKzlUgq1sFCZsUGvDaB1DKBYLwcFA9IRqzwNVS6uSZoL
xSRjK6YLD4HAWZo15Utxzub7PintbsXKXki4TKzYgs3mZ4DpQcnn0HyEtstz
W80pqXXHl4V4OHplQRDLU2kmqyavVOr/xiC+EAKNLHCQenPce1FvMtLRrPvw
Nhv18IqwYEYrDpm2Vph2YrTSAAtannWPS/oIQ4dhwX6UBa6tb0sz+nTIehC0
ny+Xa9UDZjG4AyLkqBUwV0293Eo05nNqcmnegS89D/Rp85pTsRYt1yoXOXPA
Tb+tAeja7G/2gIcWM+mQYTfSVC0GTiJLQ+T91XrarEbN2yaHglnh5hl+Hu7R
L4z3hLrHL+Vy3eLCViVGClCA6HFyceOaj+yUC+xVb//fADatMrrAnimIEvss
kStk6pDagMFJtzeeXznyp6viwGIBublDFvcytSYzevp5faFbadOuIw0tvJig
pEp6k6Uf/OPLpm17Ttk7gECU731Tmw3e8s/Ll7CarbuNmTvflifu22WCsurL
+ZmvnOGBz07+Hub6hJTVns8kXHCJMuiHMSeubOATnvhm5JRBeSlCzZeoHN5U
VmxuvRg25pW3L06UBgJmU6fzluJqq7EnlM7n6MvGXingS3yvN4NOAjH/Z5Dh
qog5qeR/qhQ68qSCEIY/G5bhS42Uaj1ZRx7kLpW0yZZCQvbRYaWOyOinyzSr
YuocBN9KZQDuOPKXDEcOE8ZQ89wWOriy4PmRGd+KxDiDSNeRrLMWeajqY04r
umSZy1mbyYvckGnLT5ufdwMkYXk5zNRJgKGcGP6hflUqJvhFyUjmC8ZlkejL
ULtW7zR0XQYN3Orqb/qwxsAsCAClPoV2KoPorTMlDwge1z2NSQpjN087+xk9
K6ZxhEj14EVylipoJ22K12Tv2VB3I4q3K987R6N3EfGWWWAHdS5a+iFJUbgg
+xUIyLT1twwxBfmskayHdhVjFf2ZoMXFfOjxpln0mbMeXHYUD2JZeqXmqY5Q
aV9raBGUy0Sf7KbtA8b/4LGtgumaRu6+Q4grDzqa7Wm2/428fXrLjO51pq76
kxQRIpx/j20KEVFy8OpvHJ2B7TONR9d6VOBe0FpIgAaKeV8diWYiyN5iDIjy
eWisRz+1+Cu25iTl/0Ud/LG6lGvMapSvoswp2lcSnHWBiCpd3wJHzwO99Tlq
JMc9TqSeaheWGn9b/8rZLk7fm+zaM3W9yvB149DSCfiRROjInJIEU/eXmV/t
GmBw98cvokQFbya12cQ1oxqRnuj8N0CPRqQvfu4F0FqEC9M5mYzPEpSeFWrI
G6sBHrBauA436gWJBxCdeXIDa2hS2UMQ2zgC2SB3YiY75sLl8GY4+9jG6JHi
vJ8mSAaXQsKMGE5B6iahmISRKDPjM7PrKGD/oajfyGZsHEgPU+DWxpcTxpIq
SGgrTdA0feUYAygrw7IXHqGjcEKbleDzE8JPOu8kY2ygUAiDrZp0ZLuFCQfv
2J633RMwxGLvXEgnEm56y36Zq+G2dfmoUA5z5OqaEHG5jpjqKwvGwnE4OSZo
E9Nla3zLz69poZJ0Rl4QsU34ZDfvx7wlnOPenWI7UXX11LIXxWpKO9QM2pOR
dEZjLfZZk9nHjdaAYLrU3rVeKmlCBc5dLXrGLI0o5p5jqmWS3JOUhzrz36m2
z/mnJSKxr2XlYS9qD95woLZnJKNcLHtTgljjPEN2E6X/3RhzX9QBLk/uC0Os
15Al5hBd4Lgmb9gAUiAleFW9VDIkWWOvuHuMcer8/E3juyQlx5Dp9agVCMX6
ssQTayxai+Z7ArGEekwy4GJlFKeslGWnKbMp97RbC0l79z+PKWA0T7j+nr8G
PjXDEHF5vqTauGw2sTp5a3u563lGfZPzhVqy0Z0c0hk6D9xKqUC/mm5mhoco
XyfyQNbmB/7sCd76Qyaac3EHE1xJ3q8k7srdk2L/ajIIc1dp1MPfVyGXf4DV
ESX+3wDlPX0B3BXDY62CDdr/dzOKGWR0VAl+qNbSZzFlk4R8fQZNTDGBw+iX
+v2jLJLUlVbpsOVr+BMOFsb1UI/LCWU3VNGeq0WjJ5Q2C+JjSoFFOjJhWz9n
Hz6lwBuXiJBblBr/ZBFFAqRyMh/iAKg5uUwjZnE7ho7QXSaw1l9oyg/FGj1P
4Okocs6j3IjH/wjVqhk77YCVQ7Hz4vsYxyHhhos15HLRgvQpjVSeQicL87qt
FkIJ+/MN0pld0y0P+To723gCYfZYyWru1Jz3mjz4IKHawDnKV8lm6qPOE3sX
9UuuNOCM8/3Y4TWUyGRGW1d0dJgK3srfIs2W4A42XXHhAtvquLQ24AVRgaoc
b6dp7CUziZtjVe5BAPjLBtptvIyzahgcow/4lC3L/qqxgeQSdsNClnCWPkR8
pOKYNmTZTMFcSQ1RyBN8dyqPIcybdEoN/aWDtZV1v/YxB8etk1K2ahy/RNm8
zFrTe9BzRQBlgt8qmpce0cckdYlPqECq3+r880RnDuKWtx1n4RXe4Msjj7ef
Q7PV9d+Bo1mRxCfQzslwIlYOQFbc3RFKuJQoJl2oW0IR6W6wC7qAVmRcDTyx
eRjRRzA88Uhut9HI7SKpb8o5LAQ9pMuhz27AW8CRTK6GDPt3dXrrBs014c8l
bP65/S7rCYU+vidRiPwHoY+blI53uSzmk4uvGwPaT0voM0TWwBlGis7TP2mY
1hCWoLZPYN35yusyz/uABK3bMQdgtKAWnDla9Z7R9sWOZDXaP4dWtbn02rWv
r8uw9A96rAoXfSZt97TgszsXJXxPPrqr8ozUqua2HwMLeuPYD5IiYg7UwyR9
YjxmKIOBJ4kqTQXCILvopxMe54zhvNfK1X1vdo/FkgATPb1x2y7ctpRVrsVF
u6ahLlGlaBoHDVkj/V8URohJtqWufo5SNm63m8/2EXdTqvMHJEDbN1kBi89y
9eKkCz2WVMzrVFlV3eeU3+CLXFiovrLfoSWN8H540TybfjDAm5LErZyBlxpB
Lm6x6oDc+COe8B0OrHSijNK8hK6snma0RiJKAmFmkEx1Cz+cUqFXMssp4gxN
vy5zT3Yz/LPoSUFkqGejjSuXfh79dbb9ILc18QbaVQRCemeLeBNT/bU2ESmz
9JF+iXpfZbv4T9h4w5ZaFbb15PQc0ig7KaTPQN7cf1eExge/sAKQXsO9DEvl
JVGkReEAVo1jTeByaCghsBcxMhLcHp821wCMnayvFr9PBvr2MbV2Q2YcfK0N
WMsk9Bf9EH5BUVA7c1HSDgZJy1Iqa8y6lU9Xr7OqufWv5KEk2syPI0mPzULs
ChUnfHngXIgC0UOhwZxNTqoJn4VuzmXnILSz7LZFA2Pl6LNkrCfYa7Yrw1Bs
ONnhtCLzsiOg/oEZwMosTgVAdEeotDkPxKKReLsJIDUPCsuC3BNFKXqYZf2N
pSXBTsDBbaM3EEnjsFjUz2k/5FC7DOmM5MuKHxJcgAh1GXQ4swWp5xZKKY8n
yjGH7SEagVPMWXjFbqYmoCQaDMILJzdw37rzbOGRoyw0wVdB7zjnX0XgZxrs
eobLrogxhYbrRliC356mRvhZC/j+D+wxbD8lKLiGTj7kJAvI3w7cVLTY2qlF
zUJNDbWrWq5eK+ouFtA34j3sFP+UR+xcsxuV0pCA/w38H2/bmvNrb/V9q5a7
uvqA6E9nZ2PSMa8ZPGTEs/vxtOhlh0T5cvCpEOtHQ5zeAXSWzh6rDELc4MSJ
xq9jjChhzBwJ+7BvXKSIWA3Lc1W49ikl+lny76Iaz6bSpH6xGTEEc/dlAr15
PUnPhqq68S7AUECMUGULbe4J2vHJmQA7+XzWi4qHwUUymr4eFqCrsJekbBgQ
cJhgtoblii1mZXHetcLbi7wkiFshtMRBI3/HpfbZ7BXEKyyVGJkhVu+gSd/S
T5M2ybIduQ/9eWWwnYEfIPsZoxL1QazXwk5osbAdyG7Z/lfhsYelcE1zYArL
aMEpzpgSvgYCLG9XSJKaiEJRtzk0Em4M9WWBqMNAouNgpLUCG5kJ+139ZqUg
8Qzi15LkRrCLimqXdXkPmA0QytEdZOlaiD1a2L0gNQJno24KgD7p0J5XWEmJ
anelM09QNFpkxS/BQr8KwSg120xzPP0Rild5vZJ5rcxQZYZp+HwcApO3pYwA
lIhNKXnCEsqWbRd8ale1TyB7psgqC4QQZiI1H/OW/Hzgljh89urBzZdBFtD0
Lm/zUvUwnvFXbIYmFi+6tyEdSliuBXWp8VAMISYy2lP7GfxMzv1L13FE3KjO
RNPRQ+aCoHOnR87ialLK+W4YCbsLYohK/yslt1COUMW6gaV+S7gtgBEnKxIs
OssKxIWObk1s8KX6tm6BKMXLps/UFd1sCZPjgZkaWTFThnZ8zYJy6bhOqaEB
lo9sAtYDXHMWOn6/x+Z4l4trCfIOmNjsHreYyW0LIlygN8u7NXmGvdez9hoe
sR96tMF8/Nu1BFt4V9/fe2gvfdGg8WaLZiRoz+fkEn2U+USs2emSpBpkjbN8
ipZ8+wrQgctKPQ/eFlqW/Pc0aCFazHP52zF6aHd3zBt8KiUMhgh/uX5kif/L
CQ6gA6qOSYL/E+zZ1frmJxTnO4wNYqQ5VfvIR973Whtpm/kOa9DLHEYXCjIr
oMWaYUC96hTeAGDeld9E5A1Y5gk4CThOgV/5fonMYNMPH5NPF6eti8LYuaVY
ePtCHl63IzKoyInRYcmBF8/Wvi7Khr1MKAUTug67P6vCRzdfROSNpSJhkamL
YBKSBbsiFZsQXsUODFZvqGec//aE/oqktiBcEvDFVLeLIMWVMQoo8790uH9B
TSmCiJZw0rqihvSK15a7k/7mfBE7U32fCgUe3WMLYoldylBbgbeTkbduzaQC
eKVUicWCuAt+dA9PEhmrJhBQ26Vo1DFBs2yo4hWOxMm6ixAFJAvnTNuIRGmn
nyfa2R58EfxzRfq4NTtvDgmVJ7VIEhFkl22vZVRAEQObWUFNYvAnUXuV46LG
aZvTIzs17Mhy74KyPbbwQpOd2j55uUbKrsMqR2QjCw7Pe9xAgOzZBHQc3X/J
ZPTYg5pTd0LGjQjCei8/kkHKQZzO5YNGz8au5eu/cur3mLnjPihe9jW7kES6
cE4MqiUlQ9UHDxGUkUWviv/+hc/cegsjnwW38TPlTwhpcvLJtfcIeNXRQnQc
xCTLhNR0IQmJFPzGHOAlbTGcjlEOzwT5Cb8h+g3BZDRsqA2301G1R2hhJuYk
9+2M4vgi0NpDh3N9zA1UjHIomvQIrNv+MnHZ9+9r0SB69LJo2l7c8DD8jJ9O
tdlwfXbGzNQM7A1EduR61Wi1yCAEfvmeTm5mCl3OpdDeZIIB8WH2zvKYXdwI
Om273WyKC4gpte98Ih6lCCPmbqVbkClXBnXUTzCPQtFiimYRbbw0kJeAZjTd
JmAk7UfZdjKg8Kv8JcWIpOtw1DZgNssYOFZmtOHqp5yExbFjcLHTg8m6vibh
saSXnxTpF7kLYOrueXIksmabRcVfUMfB/Okjle3MThZ4X5gAr5z0uBy+tlse
0qOaDfKAJ5xEPeaL6Zr1aM6S40A/7tuLjZp8krwo2uQlKK62+oDEEVvMNVjh
JfOW+Yk4mbQR2sFusXW4DsrZIpQghyb0fsuEwM6hGRgJ9i0zMGyXXJ4/LB06
KYBSkpMyM0JwuM5AIbDJSCBgtVVBNByE6YRvTSA53BFfQhQmQOe93ruP5/zx
mDfNS1ta1sp3lUB2Myv6K00RDoVJ2/1AzaPkbMnnYdZSksL5jMPw5GoLt8RA
TBH7fPOYzTqIa06yopH/pjU9ef3ucAbi5Kma3auUMDejp6sDJ5rOqIipjNjQ
9JKUCuermh3m5K2jlf/CbXjmfHnwF0mvN+NbFowT2/HU+M6tmIJWdHD/NuaH
YcNHEjCDG04gAA6qjLkdImkdTkgjc7QiI+l+nDxX+tlu+gmPbGtRSRazeIlR
6XUxq7LlZqHZ+BFJbGzADt5/R4GbhPPec25pDiMTDH6RE/jRbapEC/RWDnBc
bxShpwWtCrg6K4J2XaYY2k0OhCHcYK2pyW4VrxhIhdXzv1l+idd7nrYUkpRQ
4BW3kt2enfiKpy/e06X+1GNVaPReAUgq0zQ8RxEHCRQ0VkOFFO6mJhu1g5g6
nV18LwmnxNIdwsDboraX9L+Ocgu7YTo16ODAMjsdTjAsy5bQLDKrhd3pvhA4
uGdmnIKH5OpiuKLxGNT8V0NYdiUkiO4w758dTAge8m7FEgvRd8zDAVkZWToN
pLcqJquDk1SdrFhh4MAocpb1h1w8HvxE4L7TMx33qBZAHoXdKY9rlXX+75cQ
dp6RWzjU79Xa9cb7Wv8vzF7qkZq9JdATpm32o75FhjR5Mvlgdv5KwtG42Nkv
i05wJx6WXUh/lVzicggVv1qOWNiG0cWu/cXTXkyN1SJhbG0gZPjM9m1voYta
0bjCop3wAiwTTCDUet1tW5nMq36u58DdW6cMrUNaVWcqBFWaY9KL8/uVCkTA
QSFvP6nx00O4J3tnlftDvLRXtzV9Ct7KAgkWXp1hDHjXYg5h5kOBgeTujVmF
dUto0Q8jolrOuhvhROAE18gHrSSjwULwfLkKIyb5NysIwWGaBMmOQ2Fu2iGg
ENoUe9X5yj8kFMqvIPSJ6sOHGA12YEUffY7MVXn2ofwm271Ilq0iknaYRC+S
8zAYpZwptyaN/iY1LOxyueVOldhFg+pr/FTKNiUbPFp+lYoWV9k6Bcktm+hj
cgwoHD5xnz8T8wlBPVRzKz0+tdaB7cQr+tzOitXHoIh7VH2KkxexcC4E0CxH
bLX+vMr8mEZxaqGxf1L1o7VeuYPt3iTyFCoJgCZ4RbmvMt1C7L0bsRgh4iBr
3yZMYy0t6Wui+WTrm6WbaW8GpBf2gilqnlcFVn8MGLU5rQplPd39V1YBfeaj
ZrbRLZO5JIXyIugE5KhkD1+OGD5bWPBA+HqUDIPVxFIQ9y3RPjhF1R9PmJY/
dnENR/v9auB4hnDfj8gp18mzChvSRLZvoMCRLeoohePxaa4dJ77QsKEhxALv
JyYPFLdPJbyhIkZ22cmOPaiTVWLv+OAFVmhph4daTxmig9/MO4bwcxZXZ3QM
fq3JhO722Eru8KbkdqwW6wy+zoVdeSKxWIjleYUEUj0Q/u6ujCMnQ5slwq+n
pXOU0YtKNALcUr1/tsIAA2WAG20kSughciki6R88gcs5hk+qPIHkFD93deJT
QYJgc8l7BnU8gFXRDkRJdDFgG8ZGfTAAYKmqE3lLFj0PkbrbKtqVikR0Pi46
gNwMP3whnCOqdYcM+jKpJJxgOUTUlzGCSwgq+yrea1yy6yFZJJNiFGTP8X+q
TPqrjc6L5sZqFTC6vcE7rZu0MqLUkA/9YOqY6aA0GkmkLzfNodSHuYOftmGm
0nFk5y7FuLUt3H2On18GdlgheNUk7+8wiKHjdyHN9v64dZPzHx5yMXRi9t+w
UCxtWlrbA9L4RYep5cvPgvdetUQSeyTC0LlRPE6ZEDBiCj6HFuXF01LAWHeG
JLzjKSOjRGKa16XTTLAJxLXpMLpUkO26cnDz3U9cIOcU3yd8N/Xo+LdaacLQ
cEvItWK6VTcAP+J34E8DuMje1wsttbFa2UgB/Dmpt6T4ZPwfD56uHs/y03Lg
FUlNVWb2gqylomk9JmbnUeaAhVU3ZQEpF2QuBioTa9aHTgnk6ZpsT6Mi5FYK
AgiySS3+gDUpTgqs6HRavYFM7ezReG8tlIwNob8KU9P63xwm7CYZgpxFOqyn
zKj9AYcW5I6bKYzaff0FyGNOIMFWLW0SLERmNUENzXG5fEwBhRng6HWD/8yS
l6D0GtNL91UVnQlvE5SBBcDH/N5oOnSY6y4cTTA2SvAjV/R3C/OgU3kZwbOx
QifbCK+7C/ABzTyhNRwOJD+3aVw3hPQArHF3f8ZkpdVxlQvPRFqYW1vTFaFs
xTUbkZUciQ05alWXmd4X5tNxQ1m1DQSuE0BZ8t0ut8ksh9Jr7HYzhMWE6mBN
CL3hsV5TMEUaz/2UMB75odOYUtZK1wFUIGHIxbkNh8zEcBVLLeOnPU8i8xj8
yhUnNqp4w7QfywoHdFiz+Zsx5asyzHgW3gM9o9Uf2nIHolAHw4sEyOjpj7+h
hwN53YDV46I4xGhRgE8qI1xaUFHpf84rIHM0cyeAGTCpb9keC4xL0j8L67Np
RGP7FjggYYKvzMTnkbu9w17EPjk9SCk2NYqgVkE3nApvRxgkel3eoAmm2tjt
kaOtQCBt/DQWggGIymMCpJL4NFa2S4n0RzUTvG7vTBTcd7D6x0pDApiycRfN
WfiXOIlMfJ2gbMBQgL9zsG32YwZUhclBhL4kJ1OhLAPlBsljx91NWB9cJ2ce
TvB34opQOs1i7AFx8VEkenDcR/2K7+yCxxU7kTzpomPrWG+bdoFFxvAu7W0n
vGS0ofGdmnBjdlunqGh4VeLiQD0DUo6ti7caqihUQK+RI/CIQ5eNGikLWrhF
WjjEYEbRI29UQWT1NyiEZQN6UqoEJKdLP3Zt831h+RVc/Sb6N2eRz+RiDMHL
t6gSNyNVq1a39qkNbi5pHKdkFPFii3qGwXmsNubq+WJM7SbdKkMz6cfazzNY
WweV+sHJuqMOmZDSnRXgp90aaxZ7dzzpBV2jT5zZKxYf8Klz2RFeReMqEu5D
GY2CTa3KEaVcMW0dF4ymTlJGS2mAoZVQrwI93/hGQssDxS7kfNCqiNng0UAe
O3eS0PmGFBwKii1GbxOqsToNB264DVa6RlX9WsxX+begN2Ha7o3sid/iRsyX
MCrQ7iuRnu2YcD2nNcT46KPmR5CGNR+bMfHAyIpd8gd7j3d2BjMdxUn8XZgN
fWPgJQAsLG0MeDEXYaJB/6V1tLWNg1IRbuxNJmZebydi1t4h2vDGrSh8ZOdg
v82QkxEQzg+NQopM4QSh7ek4AfFZhLqoS4eJn9EdNR9PY3GjMAK5c81CzktI
Ae4e/5UUB7qioZgTFUPAnhLEbuEgYkItV7o5MnUdGP7AnMz/nW5324oiq2Lt
JxskrhrR4Fio5gT4uG4GrZzTDK99DCkRAyfYBmLQeqzbUMjuJaXcpbRd0VBP
drOOfu5ndoHURj4SQUhMCH6IFx7606zpUzUBxwTnK58hEfmXPhNbmj88KbSx
2eT9FY7TMZDPb2sW/C0OfnL09Ty8uDuPwcPEduqSAxwPRoGpOB0Ml2/rFqax
DyYbnSkTpIMWFrCgrQomn35cKJ+g/uYHbSUkPRe1rmB0aWZw1oK9fc/0Uo9q
hkrbM0piVGlUJjauWusTm3diwqj0BZfbLkYUpl52nsvD1LRWYwrf5G0Dxbid
KDon3sEr1+rMxWMqZBC7Cj9EJn+V/R72NeVHsjpQ/heOGk3Ani+q2cUJf2MO
DaPpyAdntQmAZT8XhtZ5gKBjNY0twd6vCLnKibbgwSJe08xBlgIelCyu/mFQ
jKnTem6po3j6LbBKxkAgi3QNTYFMfR5ieCzNv/j3hI3DjdFL0O5y9kiYhG6F
8AQByG8BdcR8dSnHwvFLOYXk/mTqjEdzEuDscKTflFM0kBJU98BG6c188MoH
if8GBik4WNsMDDRacJw9ceg9cm2rSc5cIZw9gz6iQE1gNtitmxh2AlIbsK0S
jefajlwrOxqO0apC5/LXe58xrOGYOcSt9akkTij/WNGSQgjbUQ7xmaLJLqZX
C5v1klANhCQY+2xNAOKlw5a8CfMrMjEcSgwBG/HnomjxCUU6LHfTnvQUnBaf
TULUd+Sf534dUdS5GY3URXo5WUEeIo9JWb28yaPrbR8ac4tQi9D/H/PAgRXd
Eu/oOIEG0R/2drqRV9bX70se4iMV1uwQtHNHU/WgGYcCq9hN20sg/Pkn/XaF
kDF6RKmQw9Yx5KA+pYcAI8MqSkb30+7kaVvjx4LdD8LQFy7auDzs3OmmMy8g
LmtmfcMvccPX0sqf4jy3I896PftavKcophpThGcRVT8WuLeZjCa2BXLx93iK
gRVZGNDOgsFRNLZ0gyR59KbgseXc0r8pTvY+GeAu2Z5Zs6UgbyFni/7BoQin
uf3zu+BHdb9Lo3G/fEzMLHrcUy610papQ5U/jlXTQjQypiePyDm8SQAycS/I
ViwOY+kUNPdsE0ZHUY4XEMWe+b2LlRXI1GeIiDTw+kB04yqbjcgu0GaD0ELM
Kc4O+hY+zVJsl81Nwt9kx4LB6Nm1JsnF0xlWcYWWxNN0aHU0PAcyni5AkgUS
4WhpEEXXAIsgTthwlNm7PWePK0C7w80JeTX+qltIr/l13yb31CNR2fBka8+c
9LqAtJFB+sAH4cUmIslSgSVzs4qQjcNZ4xLFCclUW9+q5f0ANQtPkmAtwLDr
ASkb4j/ndWJQTajJSKLLBEtkP4+UqDSkf1R2re3A28wb9zZCAxU73YJVlFhG
gZkd2Bj78vS+OBa+rWYsLUt2rEB7Po5fYHoNMaQm+4Fhe/B91vWOomWWA2Aw
gLwryQFcBRu663aq0Lp9eYFPBvI5qlzckeyAff6h1ELfHTX5DtmdO8RG556j
AhcE9CgJxPVbbyuUmg7DfJcqe+lp71/Y5O4up/HSVCmy31bdt81S01F0npho
cvVPURl+FAIqqA8WsGFWJB0PQWydhONt22ATGTJ9m+pSD3BBx9Z2jXBdl6Uq
RJgIP80DTUrNcuNLPKj5LZ0mRP0/4AY69Y2cwWiH0Jw97wFfaRFqZ3bFkZUJ
81Hovt6WWNGgo0+1gzaJOz54h087n0hNt1AkDDzxrXDnBS8LS2IjB+Z8SwBc
/2679G1y2D9jz+FrH3FGwIk/vxeBcNeY3gAavl8xXs/9rpOA92B9Z4hLZ7xo
x8TAtt5a8mrN+L59hY9AHm9Nv+w01m6m6bA0OpCCVX9G+gYR6kN2GKq2IBEp
V2EWbUfXsWKMdaVog3qxYs/N6I+IBjVb6btZthX1KJppQ/oi4os8Y7DDlpbK
NzRErFR0c/sncjKuKX9Q2qFxUIAcQ46NJxYPq2tgdRzGcQXzDFToJlFgW1rW
9NLIorHcDV7rDhbSWTF19wC3bQMTSOI+akvXiaNpx6eEvMVejDwIntY9wVjT
5Rw9uZJMylXhw9JMYydSmZVbyspDFB7cm/d996tk/mAYhhbgOkZJH6rDnUcc
+xwKF8qM4dRHR8T9swqgoTJhd08bsp7dLX6uv7IvCy83IN6lrgQO9+Q8UBKz
nFyyOyBW2p5RxEwcfvHEUgs5PoFVgX0htN334x9qB7c9+o9imGrTxuANgraI
5jvV9g3UQVFzlUj2zS0u81SIOWVl6bNnUWPhP5wFhqFeGaT4ex54qx5kemic
Z+/pzBBSJhizXWRfC/UBQkMAucomA4HIEHvgJ1adusxvhscsR2/DBmP87ZwF
S6c4cgiXTaLc0ErvVQmlbKh3fgg2SyIxEjdgDTwZW0pq5PXoE/H/8qmmLZBl
GXqUDjTKsLKtWte3BPP8msq2kgH7P84MmkDe1yH3OMwzeSriX841NRPuc11Z
y+DCNSe/tvf1rMFjPDpAym4NPcUArR03Eox4wFx/oft7ScEefrXnSPgg73ra
MlQxwo+rOWmfeMvh93vPyT2MV2Ky9sBmohNKLPIi0ZVnOEVMh8gdLi5e3c03
B1zJbnGeEH2tHbmrcJq6/Nu1JSpMfOwX3vFS2+VgdBKYPiDTzZ3zuZ6IuDhr
Xg1xHRSneVGdqUaRiMLdhX6OlzJtX/l4uEOEMpSIwsW+cid1E6LJvBbH8+JF
PGn0m/sIfRK7tDXXxlJOXaFHxGk5eijTCI8EwIdzyMRlRgwNlXRko4Xc1Wu1
vVEReEmu5LDG6SlDKc6BXxVN19HP5lrd4ujCj+Tv/+nUyBKlHA1APy5cBy5N
ymnDwy7M3lN0AR834JJorj9Bu6Oi19iIiCP8zaicgs1TOvnvsZGfAdV906tC
o8XTTIyl6lxvRLiLiWtz6Z8e0WV60SR9X7stA0fsROgeI+fXHZh/E67RvxpU
KeFVnmC3XTVJ9MqfLZ5PxMaWKv8spjJhnnB9yU8uMzX4q3VzyU+BpTrSOykI
TsfD+3DIrak3dKf3SO2SaPkVZcsykszrYf40+P5UEV6owLkiH7rUYYhv0ept
nyBidpvm1onb/UUlblNZxjoOyO21m0X7/quhLJ5fB84pvJ7pzYmcqwwxTuj/
Kldc8oEafe9sTI1N43pBtG57N55fTwIcLo2ocWlJvNwndx/0Xs0Cc3LUPDeN
C0FefPt/BpoPyrFFzSL+FdnC7S5+1yWCrCtKE21DGaCddWe9nBoHdTJcOtiR
Lc4Ki/Pe5Ky/f05VV+FsWhxaWEEzGoT70EjmxR7fMjH74Eiwjj601+Fb/uTp
IdHneDF/7ql2dVkjpw4bhfG0RurdyfhWmDskvSRcfhzDL4pUGjEyb3WsWE5L
zkpJOQJi75t2SKChd3rzg3KsuvfNuJwQjBuCiOh6pG7Ri5KxcFgaveSvzBJi
GA1mqzWMoMURjIHq72Jg06LTVhmnJo9lMMhwc45s2o7jyInrS+bMsJPh8mYd
M4pjkzMoZhN6ZvgOpt6quFOcQUidpJvv+S5lHE5/w/uJCfLO5EJclywMOMEx
IyygJJfMnzLBdQ2HaQjjnlw0ibIMWsq9XJafkoHygg184mTUfaQHmoKtgqxT
bp1jlLb6Dg/usOyjm+ky7kqiALdZwU5wwGlDy1VjtYu7CFnBVYUQtnHZ81oL
vNItxJXKbHfAmg+CLvKLz5JsGrkgdFqYwQoWF6c7Zv1Z1VZ0KI8IB+rUpD3l
VcenHMf/aulT1M9+lSqxAhwcNKtPushF62n5j61esajlCUSjMyZPtBlJNh3n
ZjSxElh1VtIQg7RdDKgw+EcTsSpW4SPIRMElVhci8BTcxm9wZ7OJMPdov8e9
C20yOYDWyvdeX5F26CRLIAR60RaiXEkSTL+3ElIPuMuqtYvkM9Eg/FkMuwF0
mN/ei8EXTt2EtU63SSNPp4ESiyYHLIB6LwPEqoMFDWAGGVapmfBDU5mVvbXF
MsgBs32VNhLsCUoikGXcE97wVmnrE9u1kWQbnkoXwJUE840EU9wBOxjZf8b9
BSAniQfN0UtNIPucmSKu8yD27oY126xKCoZ27VNN7y7noIoZUpduL4pcseRk
SKQeiPa89AXlWk+4NVGUU8n1yJdAsdH79CSBHxFYTeddl/4UYhR5cmx1xN5D
0lVnKX2dfeEAeQBp2Pp9Yn8oeAECBgQhDfNspB/3lR6nW71Mfgy6o0yfe8++
zjQ2phOyejR7QEbdZg4LlFei0P6n2IV2ym8tuSD+wyVwyesMe19Odm/x2TOp
Q5MGir0yggo9TkMSIUNgPE6VCBXrqeupomkfCiE9njLHDhhhfPMEfTjKEf00
a5/aPvhLVJEZ5dbgiAvTUpT5kyqddEjntVwJT+JrTjx1XuGvjrMbFOSvY6d6
IcMyS1nLlFx4DJmja380i3VykRuJcAPVk4umDytaN6KPldgpZXKN0AVZK07i
V+cMT2Ghv++5M1T5xqMNbSlhWKFYltWR0nU2rC/7WWrIED2/baELEU6QpB6I
kwjCh1k2oFjcZIfjofMSqwyx67BgNZE/owFNwGpEl18T4G83RUbMZY2tcmCy
TU/jmAPs5XoHAgAc6U0JuAYm8obY/lam7E6fDPQOiyWKpbTxr9hkECMznmE6
KI4xqVNo4jWEK0ZKHhM2hz6FBl7G86IT1hQP5+mYDDzd5C//e/dwPINDbf+0
276TASX4r4QL2+6+a+lAkYlMF6LnSj92MmDpsWexmlm8TLv1dVRdlhkfIgxo
+p/WJWy9HLAkt8jT/89pM+4o7BS1jgecaAhlAt2ypVlDh5Y1/tF/UEBQD54m
DsKeINiZDkMT71j7exUpZOcHCrbp8pvevhvQNkZO8EPtfoGfZWXw3XwRmS4r
5NnSnCh0HIoMmgiPkm2eMYIfx1rBP4bXdN3gjBVICjqftJXFAWMJbRAZa3Bo
Ek1uFiZtC3jYjqGZY4drueyGqdlCdyO4goIBC+eEjtUIRckR7wQ1wCh0Uuaj
eJ90PRvE5gjdBruoumu/wKbQ1EPvTPguFCoeQ/j9IlUmjUEXQKyKsqwyqV4X
ec7EYf3Xak3eZpov04BTv1nS+YzKta8YwLqHENKo8BDMj2g25ZdUaqoIm2dr
sIS8jHwZatSgTO2DYr+ZgeInkF5ua5oWpfQKGGToG7g5DweuxN8AWAQL13+p
G9nz6R+BszyohuYk9W6toS+uclRxr9zMs9J7gXMOPuPYJASh5/KPWAcNZwqL
gx8s+2XfI9msbK6NFRRDvN8SZRYP4zL3I53A45n5+RjHnu/jx57PodaZ/qlq
xeMRATgjdL7OBGh5bSIWU0ysAnST/Mt5tYhWFr0p69vfPkWpd2c4KA92pEe5
rZbw0RBl+vbqDgV7XJVS9XjE1ebkAa5KoSkcSAtdidjRuZpEn1DudLSu+1k6
WMGKBk07U3uaeWRXZvicW6fUa4gZSwDRlBgEusNQBnszcn0GW7gCFoaGALSD
KR/6m4tzp1wYNUwYQcaw9VlPg7jadLxPzdT/WPTK6pOxJ3YQNQil79CLVlEu
PchQ3YW63oBvq7Tr/Qp1LoFsU+QihSsGLVjuF9sCycH0Rpf+ID3g31roRFx7
zaln+yNHP1yVCzEIneBLZecw8zX0TPkzQJYt++GNnP6i+6NyFEiOg8ZtSw6l
kKkZppIyUuGhMmEUK85N/9prAUgiNrAPLWloHy71nsFvJHa/jDoaY8gioDtw
XfoXvPMJ1isVf6GDsmW8I4JGT6AUEolBsB90k7Cn0Xs8VjKEH3DsYldcdH6C
xCUosJqOWIyw5j/51LvG5bzti0My2h6WBX/gzmhWIDKdQL+BJMVN5ttid2Qx
SUtwM2YRdO9afdfx8duh1D9+uLxRoI/xL7re5JWrQVgltsceRkUtBRgClTyS
kt/M5F+4EiSmqSaqRDkhMpiGUPEQM4SAakLxH1x2YvHoQOMhgqK8k+Q4eLhB
dpjzTAjQJl5Tf9y58FXfmPlIabMBys5IqOqS7rnxxgqO4KoXGX5uLBXQxxMu
R7YtTkTlIcAFF2BAcRI8HN96NsrhSI2PqCnPMiBXyUDRP26XPNFtgCHVoQzz
4ttyu401diwI7KTf4HB58uFeVtz6Cppq9icf5YdUF6maJ/tfDH2roRN+8a1Q
T09AcD+mVHcDmW0mrU4Cbo+LXFFapp8aXPlGKBH53TGcXgd7yItdCk2LdRgu
FhoP1Lu/ZoMd0rbvnjmzv+ep7sw9Afwn1Ql6jc7qaSFmJLtZCXQ4skRbJ7LZ
I/PRVJoRULC3V+JL+ukGs8RKPFM1nmUIMWyv8zA3wghFUex1QCPRn/I7yyQa
Sv8dDj3CkG1x/ie0g32kwasHLky/dGI6VBanMHd38zuCk7ubGaWMWVMpmbUy
iE594plvKvk1fmvxJcYEvVbuZsUcARuRwdSPR7hhkCuRqz3uvVyq+ytLhxQB
EsA+PDRKBmeWKeaOQU4pl8gKzSpQViDUCFkcStYCyDArr6wVg89Avy809F84
PD0BzyPMp551Cqd6H7gt5+mopJ+y8gfw0uasLJLnXT1P/HRk1XAQHXfXUzyb
PRg5JWqIfA/u+RQzzsIFe7VwJVpdGkVJSmmzoUngblHZ9O+yfrrIqYUjsJle
q5IJiiQq3G3dmb480spvO/jKPINHfRcOi4OlFrSBu5+ioKA2EOcnqFxnS08w
cZeIfx2JNcvEdW8A7T4sOhcXn55CMxV6w/g1ebduL/Sq9TYDIZsbRwW1xoUu
hoj6+cqVXJXniM1IPHyiNNwG6ReBappVS294ceTJVzeMqCYmQ4rc+TqSwWhK
2upC1wjkcu+wwtfy4K76ppFvwDBalylfqKr+1AqDQ3FmvAa9RPQnxU8Dv8yl
pps7iC24mpxDhs/5cPL17E7RIxJzom6kyc//t+Jjah82BBzNSzQwG9H1njDD
oIqSasq18hpsAKJ1AETgV9/CjCizBJ30Uve2hdCeEvPPh7xo+1lUlBP2VM9q
fnOwlhQe44Lcvu9neYgzMaeli71rdMVKeRDLjnF/ohMq+t+wgrnJcyS/6iIT
qC/P9iaiLTHo+VV2ewQW0WbLccoUj3Tzg9Ks5lyaHJp88fPBW8JUjzycRJQi
z1kcZtVbl5b3/FcmkpIw7MHktsphQ9LKsw6OYCE4w+SfjUC0CJkkONYivUcX
Zpab3kaneyk6cKqi8X5JYP6gG8DN9WcmQVLiNBfZeLmJtLVYgCXKlsJY02qN
DRo7q8k1N+5G2Rw+c+a4paheSjrCmBZObyt9OtLbEdCGxzrSIPz/XvLFwC9t
SFRjkzVcgnOupUtxhY/097R5mBFj3dgJx7fE5/0hs0BkLzXT+ytEBZimYtT9
BHj/UAVi+wVBTki8DvDOLLtV0BFj5UrPEQu0Gwm9HSuDsi6Gy1DaWEUczz+8
vtkAXATIA/VQfYfcWcQQzeR9XIxH4QdMlJPlx7vMbAThV4u37TL8JnXK5npg
xh2HXc8AR9uJPRs0dEsoAPpqk1ImWW89iV4W1/YFviGcQ0gQBNkDDHfpEI+O
RUopfLytGt25p/9n7LSKdd01CuypPvRbXloOpFZxSe+rq/vGqQuCHGUAXyDd
Lp9wVcnU7FIMi0Gual0HX99VA/AyCB7dFBmA5XCxETZE1PM8TidmehGeKi51
FBErecK+TGb9ABAgkZmzkpcIB9Nh2sYElN1+xDhYRoOJ31Jfm9Rx8AaVVqqo
ZIzRgRRk3gEVXteIPsQ2MyBGZlHUk7tqkeRyHsojdZPD3/bRrhK/gQ2JuFEt
CNKYHHziML40/u2sTKozwg+uq9EudLcnWdRwsow2sNflnUmF7y6wdx/tmE4X
ttMDBbssRaFVjTMEHyOc/W2FDqGxV4/2YiFfVMQA8i0YXnZULO1zE6Gw86tg
EFva+Qqsyoq8t9KXNcvAnxtfxSRAPP/87SFp87kDSmFJI6XLXye1uFSwWVN+
HKyxY76IH2bFZfH3cOq5olSn/fBhQM0uIxoKcP5zMhEZ9E1+Ru/BcF17FlaV
JCdsD6u/IyS3b0cACnM0DGKqYAHCC9LjcaTBeI7hwC2aHW2elR2HRmzpDpLX
AZOkPq9K81jzxbRKDimtwNjy90Ayj9GE9p+B/8zyNmiL/v9ar/pwMvB0oBL3
c6JsFtlBe/GMlWHUwl5equcMVnFlav3C2JPWc3zQBoNHXE/kMad8h7FkJKuO
49cHebd9t6G6jFtO00GCMadIvv7Iw4PVPfSlYON8KpLWz06u50vKHqa/tde7
20fgUYsR7iiw03by2boefdPs8zg8odRBw3vdQKDBoogHIoIPTB7RBzGccEyU
P4801nSsVh6I4nomdaSnzkGobPwP8WGmbcVy+UGn18XBkRwiw/OGr5CdbpS/
krQgrvgIs4uxNkKcY+1F+PSrzsw6ZxNkOe2gh08KX4mcqc+qfpMJbkZNjNJ2
aP5vAIKpJiEkCCGiWTzuYaSrfwQdpvpwxYAugque8yfgdW9OPwhWiXHlpTiX
AMrhYcCVLczVPrYp3cUNk3URbYVtW0rCgqZikMTUFnK3HEEVmrlYWbb9UwpS
Ka3qkjtVQ7fa3WyCIOfxGBQ5XNzCr7/QtT+0WUF35SCOxln7BHLpRCYeu5My
19ezC5vRW1/vuQbnYKFT7i0WBZLjoaexJSJjP6PTiDyr89YhTgQvG6cXyJoy
QgffDyHVwnacjgyvNLBIj3KXEJYaxpLwxDcu/xc6aW2ZGcTEYIj6p1uOdEKG
vXO5vc7QeNbqwKyPEiZtCW41Oy/G2s4FtJwMiUadulQJgmGMLVqKK3hVH+fG
jqpzZDq1WV4HW4bRQiWBbQtPCZLQJFfWhFCxTU+Cx+N2GOAG1AjhzcrgyOA5
h3HzIdeOefHfEsFuBvAoUy3JP536XSBMr2H6/8WrmspFWOiHAKp0w8KqtlbV
nuq9fr7FPJcHEp+k1ZLbLAzvoHf+n+QiqwRHYwo/TsJTy4rLh+Ane4rhCpr/
/D4LzC8JEiIPjmNWGPrEyLIhCDHj7y3sM0MzNH6zPWZWcXfsbUQ9fYs9icBc
H8Rl3NjeLMHr55JGTXiAKJyySX/2PdCtXgVjJCzZtoiT1vgbKBn167ZCrpaC
t0V7XUtxdXXs47rdMl7ytaLaUotjNFUel07J3IbSl5cKijt2ZxXOZS75IVeo
yYnKxqKJK3FidYvz6wwgqSVa+/OlnSics0C53KGbOvnz7c1ToUndMVeoA9pV
Ku6vHkBLxlri2Zoc7q6sQhf67KtX7weR502ZUlVGs/DTiSyKSTUZm9nyXgqB
Bn4CW5lpTH8Bp4OkiHSVFngU4vIkzd8qOJ7z7LVLsLcIk015FkQJ05qTyTg+
UNWypem9W3U9KR/5QL/Xm+AAFnRdAXPuFj9CHTozwAhfJdk20IKXivvMcbgr
u2YY1zX0qwewSJmxO1keVngv6tS5U5mX1GKFOAMqahfGPfO5NRDPJZxfOGTy
HdbP8n03dC7ujHCM5CwC8tw+2ZbD4JRgoeNGHajfQRfp3yp4CtIdXiOmZLPZ
mhAn3twk93oeRPbxwELZumwxxCvNxSZlvnqxQM9YGW2m1SGyBCyJ0b5WTojj
zoBAy2UCXXZyz+/WO37pgafLDGhNIPmExXGUBM8DwZyYI79kKUThZEK/922p
B63w/f01/CTsij1HsErqr4jWsp6C0ULAiyy6+tHf1iLeURcqOvjJP+X2USVw
OIKkTXJEa5p4m7ZzROIHE9c18QZCrvzF0+qQM5MEMcr497BZ73ok8XcDLspa
AFlkKzZUVSSyBfgefesuUcGEs0wpxEt49P7u3T+mAHqzRbiWtqOvkpo7BAHc
d4r0Dakh38poh0hTR1IfXu8WcmBNnpMiyPoWz8V1CTphNs5ZTuMyvEZZD6QS
woTvOGODU/4rO1HlECebLxpD4N/JBQ8IJ8zEsnHTZV9rF++QJcgn5ux0+Jlg
xeaxc7AmeLiU22mMmrqcHOP5mV8ufqdYr5D4gHyJgGRdJ1wjYyfhIkPLDZON
aCuKhjtC2Utfih20bYV8XMO0RpmkEPkzD/L5G83zPQ19SeROds6cWfi7fZGZ
H8ijxDbbgEeKTZ19r5LFl6hNvWefwGqmLSwez8B+anJFVm2K2ajeCAKPQ51x
m+rWtsgxJh3ggzo4bhUEzUuzwk78qAfETlepmdS4Ppmm5BOIdGzvyB+Q8U13
0+rpGibMBgjSxPG0poJuP2hmAHCMPUO+ZyJDHs01xoLMRUBM3l3YHa8qAYUu
f+Bj6SbSLrhTkPOcTOORV/KwdaO/MJ3tWI1UuAnj3RJBqnXZqG193ouXzU32
eWxYhLrC8Xcfi9wS6lM3BPaXZgtA+iDHy29kQmsX84FTARVhkv0vBWHNCBDb
gKanJNMHAbPJK+kl1cPNOgkUOLJPXvnNlOqkw/WQf0XQSllzNrRFxpxogavr
lm5pf8cOOb3ZaE05mIxFQhwUb1kt12umtzGfOUHUQdEzAYllO0nOh8MUJteB
14r3fmEesy5owf35yfa+iGveciEIPIUdiC2zwvs8ZPuNzYgouhZcp7r+a7Gt
P5N2tXJKvuLuOHSpdyWMk2mg2vjFhjLNdAKzEzhkBGSdv6MmGjFluWRMMgD/
4oACfzI5zPC6demM/IntcGTE4hnrJyCvEi/iwVXbzm6K9GX2NvzRjUg+QHHm
rwzMiUknx4CNcF36RQmdj/3BLO/SmJYFDd1QS0XlUU/xImJPuTQeOzEhMEx9
7Cdm2liZY38CMlpFqnkYcZd4G64GfrY6HeQu+yBlKHIbSuqDf6Z6zo++ost1
i1Tla7ddTBYhMaDoCABqPq2bAUyHPahQO3fdHqVdITsX9Fvo2W6I5AxSP+ks
7gcuxL1yONJqZzQnc7ZHoc0aCgZKXhKdYCcXRjwiOOS0Rp3eizQCZoAj/E+M
16DpXu4xD1K6da8oWbBpdADiF6BhqxkC29JxgCtQuNKRg89XNXlCbBH5dlit
MF8kLoA5OMEEPsOvlADPurRVkFicYVuqJ42CtXr44nZCxd7n8vf5EDNSU2Tc
K1n6GE+/wIIi+D1Gm9NbbovUPjh/yY9TmPBUI9cs6ObybP3m4az0A0IJhQTu
aCFyq1bj7AhykFgom2z5bqlM6Y/MXCgQgaKdrQEFe0RJP3/uxVANCMr6pAWz
eP6Rnn7BTpLAeVnXBnkH2oAAYkCYkupZrLx2NIbTVX5m8Oj20jXWw1UZSkSK
b60rMfW2mkaqkyl4sjk6dn+fUL+Nx+T8sGnGSLnFq74RSJ7sys4W5ox1jOrk
5fl39wE0eR3R90Ej1KL0d5acXnvAduXeAFHDdCHF1KaXy4Ra2YonFJHfzF23
PpzedLGZC4t6mtqYejgBBkN+n2tHTinvdZJh9IVBOJrcc3yqcpwhY+wJDRut
oIrsZGE47K0704gwCqz/5O64NCGFTeMqC1dGv3mMiH2L9gjfAermEZiQjGU1
DnjAHApW4+APa+YNfW6vbB3N7r38O4KM1p1p43uc1gdQU58ga9g2GT7yLKNE
ZA4HrKr0d0AOhv14I4DKxBrKVrxub2iYYya1k7KKg7PtohUEDSNHGeDSf+KW
s0+JopvdKJ3ctAvqEJUxrMNOl1WRwQgC17bV9JNhUL23rkrcz4THcDa9YUI4
s7kefBXQCxag7QRivgaa4AQDTbCuGDOq2I8H9GmUBrxNiAPukvXTUSv6oeOw
pWuMj0E8vLZsT0iYpB+4rMycTgkxYG+l4KXXXkX6WVZk5UGoEBl5JFlSyGtc
ZqhlNfoF4a+2pmbRGxz/ks9iDP/Mg2HgxzWLn7xFxjLRWgDOJaTnoR3PMRUn
JGZdXS8F5RzEAt/gg4khGnfL7XSIhq3FPQ6pIKnp8yGg5jFpiODUM9zBvqxc
bv4HwMjATWJGs4H1+O3oBhVBqSdOulwTyOH5lSGmYZcCA0XXoC84gsuCRdjP
KUUklQ65VUiIBhJ4dE9a0ytadJDn3Mriy7nyzrlv/NRGDfHd87nHUpisDOK/
+XfUfHExq0vcvQycEhC60nlmDe0dGIjbv6De+I6OsB7gYW1JFyxxI3Wzc+Ih
zFfJ49L6FDI8q2Ih7IQG/LXjp0v2vj/i1oUvy9ezXN+lcpHJEo9udECFdmI3
zkMMFrU+9g84yU3vw25yp96LPaw4rqNz72fhSBZDet1VvWrS8NKJBspOdshw
lkzpdxG7/xtEMJB37+DL6b4CML/KU1bf/USPwX/Cgz7FTTHmjDFXcoptOO2o
rkYaRQuoTEEHt36NXQoz/gRr688xhLQNXCK9Etv1AGSYA8B+OKYvGqUkuG3a
1fWtM7XW2mLFOtej/+imGoF+/Tf1Pw1VSiOTbhu4EYGnF/wfmuxim2BfW+o2
uJtqsEv/lxUO+ZalBNwLMhh/SRj9TOhv0vVlbw8ETf5SxapHcAyWC4SCsh+a
yofnjoiAPw0ejDNHlzk0ZUfp1K8jxYnQBRPFAZ/Exl9EbvUVVZrhYZvPlFBP
JsgEbNdhfXqo9QQclaMQGtkcvouGzJuXLpb58HoCSTkZTncx/OH97wUYZiIA
nSrhRsv6p1P51Iq9q4lIkIgnGXDNZbOyjtl136YtCcrcripyOKH083rEgGfn
cUcF9dknFcFQzsSosXrvnXazMTvXHGodnSXzT8ghfKTX9aPGaddt3LwcKNA3
PYHVWQRU2WlXEcliG8jEkrnrMJVyvPYczjnRrsoKmVIbNmn5XfwubTmVV7FF
hJO5Q6RtDvP5duiSzfS11EClcNrgfMgAaqxJHPCL7bPIGwQNaZev2Op077B8
gDuiD8MWAqXrcxkLQVf8NqQdzy/flFLEIe9P4IwQxKRMr3uhscuzKzyz9Icp
vNmEE9JTi26F8tJwgQJ0UfbqPmgb+wiDZRt0QfXJ5iuS9cCp4ep2bCIVwiE9
O8btMVjY0uxChHrvhXBV7OPAzRIrBBWKHAZTwWuowvxJ6pQ7LVNEiY4rIafA
/WcacDwEE7eezFlQVMlwIXH3qVq7vwiWRjIv/8EQw/lBizZRKLr34U5oiFyS
E1hQIA63FV34Ad6N2ki2mys4ppriZ66at+CHUJTXddOv6ORQAccbJwtcyiUK
ijaL472ifFOdrYJ3Forng3NIFpj/4f1lmIiwm4nE6qwqJa1VBJ64mYx/EwXZ
Xxa2REbDovW0rEDwtb4z2N6QxG5ZUaLEQN+68a1dQ2/ats5ZfIlN7/89MVWI
A0JoDXmG++DTTkyvFopicEmuy/To0myntKT5w3TGp8j7z9Ni9fXLe+TiAfEs
jcL1MfNCMsaRUvavcd+7fRmwHV+GLvr0SqlOInMWqAgL3qT1j6TANnvRACj7
ZAwCurSdnTWrIam29zBNn5+tVZdi/nd4+SX0hjWYlTWuHmsJcWNyzAa4/91A
XH3tROdrt0PaaVzhsycWAUi4KKQbwqs0IK5YycU8UhB+V5KC3xJSZWvKparb
IZ3THPCovBHlJuqjKpHEkdvfiIZsviaxhjZ5JeSvhnsOblQ2VCL3wuFuVQ2m
QC8a1SKxef/QqXgxRKfkveh23nA/zfqCtpHxIcBvpGLtnBFrbdosxErV7ccy
mgkJYHctNxq50ucPOs9xkXHKDwwDbumHropBOO3ONlwk9O70PaV04DqalQKg
Ly+eWeVM2/PyYrP930hbK1u+CZhDuO2ylh+upaWRf7ZX/qzsG4bnAZ9zeOvv
f/nMbNoeLur7HygQdFYn0qgqk2pilwTNjNLme0dl3nCcVZb5BminAijDzCq+
BPJL420zvRwSMM0vJkAcHGHkI7spGgrvYm8WXvNomoxp48/jTZunKn3hpkKq
w/LTyZJJWYo0gzx8wREfsV8gfQ6hQWs5kPjV12KxH/EJyxZ/lYsfZZxlwJMq
aYEIU/CXUGYpLpNvMWdRqMrQTF+pMqmo46kmfQLOSxby0RZWtDl9L7lgx/Tc
uu6gvPEpcpbk5SbIyYu23xbAJYEpBSrE7+cJBr+d6f8UFWpmVLXEG7za6/Bk
Q/5F3Da6jxw7S3bduFI9MPhpvcsp3oKVxGOUzot4l4q0QREro/Na4wCBSPzE
bK8f+D2ah/nrrbOD7m4nfPeOTAannaCM05cPM/3VRQq/T/qHJpcSY3tGvKdC
RLmVg9UNZ41inY7INcCYJhS4skG9ICT8V5MCaifblVafI36s9EIUfpgKVD2n
E15qJZI0y8q3Q96mru9bQsBOe+cqlZuSTrduz+gUNGmCDcCGd2QFTxXojeGI
tuJfCAQjos4J8+Sxl+E0HzR5jauO9toPBncef2CMfzzQy867fdUbn0hrruGK
0rWMgPPwPwnQMzRM+/6HimzFmOTAlT0Wtr/+d1u+/OAFzYBeCTJUZnciWsQZ
TFSzjobh4GkUcBdtfM23+L0N6wu0/fXCWF/UwodWU5DfJesZEtcCknqKw5ro
AwWmzVXngyqcAxUUACEacJBaFyoNnzizXXcd+pvYqRfQTc6lnkHOiMuwxQdc
M72T4YcQcfpswnjXLsCb8oHg2uGRwc0ZOdQjj4YYca/St4fNcd3sKuv0kHak
8gLspBHSkxI2XQIMe/O4PArZveGg6S0qyxaU0K7YeI5PSZpyeHrxd0z6znHP
IhlUrUb8xb+iEPgbR2rGWsURF8Im6G7WM2+IsYLWp1cSNKyiGu4BqJ8+iVJk
DqlQgOZYWJuiBLevtaQ/jF7BdT0eboKME7Z7vrN6AZYe9lTilRTcu9j0QuST
9jrdeB9EPUQuhVknCcoMMMkw7xY3fiPGFyrm6gHENt8zcRNTmZWLyRN0dO+x
TVXh+/e3fDZQj5E5yiRXPvSq6NVdaORrljlobiLtshZ+L69zR4nCxzVUOB8L
4aTk3THHx483iYa/2zdHcs1OzvP9c+VTZFYTAgHpUR7AsJfK3tPNbQctmzNf
87Ag1V+u86BBnQE4W7E1UXXVdd59oAIrNBsHhc2RROwBwvZg6QqJvUcYU5KI
Em1HzbZSSbyc0Fy/mMGOKIR8M8mkx544YNa2sTHAKjfUTcBSYNcxv5qI57qT
ajWVnw9As4UWZgliiNkiJL7w2+6wjyudMq1Md2nOd7VGDM3SW7xIctut2Fl7
6O4TsDfNIDMy0DOig/2kUuqtFJXHQR69q/d0KtxnKTy+kNY99/T41RIWMZ7s
5F5geDpQUImd2l0k+mT4QH5qDDOV7GQYB5vDPuClcmFEmpqdXLD0oGwWOlgr
9hGyETi3GbQaClcsjbTkvDcG2gcIPxNmu5HS1dQPvZb7v9btHopTiR/M1lnp
oo8HyIDmKx90gZLhas1/TGDmq0pG2jTf3RmsAOBoRWrXo0yM8gvx7QXuykEZ
v6a6hsJEODUklVXb7+odVoOnlnmMY+bEXrYrNP3UtV+FayBunkWiSOcVNZUr
ggOc2Rl85+kHml2ZmjUJfrZgUVOoR6WwIaxgM+WcdpA6UjELB62EQu1JOgE1
sbjJmgVgpIZJ0+7M+qVkkeAa8Yfo03D4KQHES5EwErZSRK5Fc3Khiz/bClsY
o/Z24rqlxSb+CyvM31HteB5QWRNThQuMEF8lkftDPk2AknRd1SrLzZ0SvNpc
irGERKaA8ZtaTqEmOK0REn70CgPsl4dZPaN4H4ttICFzKG5YdHYTDHSI0f3U
BMokJ5xbDFP5U8JHzj490SkYfBYiuiRVSeL3MVPXd5+I/6fnxxrnKi0y1hq8
JP6c8Nk39j4eFPBzexdspW/ewXSb2uwjWWN3Fvpil/Qa7LlfE8n8Q+xpTdyw
ZawsrXynqtYgiL/c8+drSGF9e/AJUqfsfhwWl9ljEWu2BTDAMTxq0Mp+43vC
gq9dCnhc+4uLG6vUYStWB0vfBgq7hLYAsRS6o24vln3aVsG6Gv5kvnFo+QX3
/zxOGI1Gq1Ag5sYKBg3//jug8QdlXjD8t+182nndwa3l58z99pOJRwWMn5cT
bEVaIM7KZR9HucQllXaMKPSxyFDakrrH/fctj5/R4Ae213Bfw0v8jwN9oRvX
jJClYnmcH4pCkw4GANukyYBJFJw6NbTOBOCtnnXQwISi1Td7ek6KgB9aAoIN
UGEdcfPuGMU6VsSZwuG7XdGYFGBM6VMP24Uya0VNi8C36KIAiGn5iFcRbk7j
cQF6T8tfWbiV16YW2ZLoic8O6OfBzHa+5qv8JmtHjPi59OM8c5ZGuu3Oj+3W
Hhqh++8IgbQEEKYCMY8KAMfJzdkbq4S9uSFIxkQ7Ql6iYtkWG7gjnuhlEBJ4
IeMRiL8i4PK14ru/YNsDaf4bs6eemhbkiFCs2ubprHCnSAfMPx1Kk60oEUZF
80ea50TZ9hYvn4bHgPnX/c8VTc69op690iTU1UrLAW69uHwMg6UVx+zBsoLW
4Y1R0Zvf8Z8FfDmZmWec/dpLoWge0MP8l46IoeybUrZrogHuOF3cOERoBaYX
4vIyZIFriQQ/IWNjogF2z6yWTWkDwjFeMYFhbe2l8bEHB1NiN/PPBP49jcu4
yZ++bw1GfbiY/PmsOLKWElIXQwiKGcIMz9Dc/egn0IZ8ACkxEl4SJqxZ7OMT
8Rt/PmFBq8NF95T1R9MXvU8KEMPmNowYteM9OF5yiqEaUIYLMGsM4Mvz6sq2
oCThO8j8o20+f8wjcPSer3pYMkrGL5VwqNvOp6GCFESf2NXgl62kceEufCLG
d6zgmAM6JSdYqlK07NzAxf38WQQ+w/upEZz2vzf4gggOqK5cZx9v1wj9Ek13
I5Tmm87RCGO/Oj3O89jopBJp29UMli9yJWmZc1qIih38U/mOFwoH7eOv3yye
2HF+e55lUC9TfzVH10hSZ7atyCAPHA23LuHQwSgpy0D7mj1jTeJcb78ilJGi
jZDsGzXrodyoUiv66Ver8mxbp4y7u+dPmFWmNSF/+LhpKdegWrH9FifuH93O
TrrxJANPrIuNCDV8y7Ka82pn5RDWnlCpCD2qB2JDxySzRG4ptKjJKqjpGAoy
WyK8AqdTt7LbgpO/EuiDP+3qQQELPo+k+UK4Ar3TzApqzGbUUEIM+30f0Y/6
nvpnR/nHhChG2fXbL/Dryfowi0EinhNVBDfUXoMrSYScsGZy+iTdlMRJTY3j
wxaMR7vP2vRTFSksARAzfUhHAffpK7yEYbD02mbgAdApBeqOg92BW+YY3qmh
3Zbp7UUjz3JoavTUqVaQtBqy9K5wMGtgSMbKanSzznRF7lT/1sIXCXawS/3o
NMT43ZPulXlcvPH/M8pz6mC4pizHZsLe2sdHSSCuXFUAoK5tU8yN3IDZu9xH
ssaACwDlqQszNBdfdXw+FkQbK6rR/VDd4EEPuHCkFDNiRdgsZ2JoanmKyAIj
nydxGo46nGy9qy4MyXVMmBP9FLObAzuNDBk8y4Y6bH4rYXxjMnrfVJ5pekwR
FuxeawynlXgLEMLquwshPOCN+Rk9PWdUv7r59aFaUgwSyV1AtyqoZRWdcfAi
TgdVf0fg3TFUMvWqXjxiLxWGqNLUxlEf5Tt8bMCfin/qCfuopI0jECE0ldh5
tTg/bsPKxwz9eavxXv9sloejZWUl4ifCI2k/Ztg9hx4hqvYEFQ91Edw87enn
pQj9MWMfUX0Bs9uETZSvd/cpLSPtJ7YXcBI+MPKYbuBo7zjIKCz1DDH4oSZE
X9umuI86LJacfY5YW/lL+QTIHIaPtr5am8vhbhXe6ozDHhgjGaoaFXPcVzRx
omauNWPjeQyHJ6uugCq1psAHG2NeSw5lmR1lAgEYBIX5ph17T1y+b9+aEEIO
AtGN3QKfky40KUzRzn/Zusn87RiLNs9CnqJkcxVY2jXRB0yy2Krk9abkyycc
Wu/mXx8i8q0z1SKXNTCSHidd3zS8AQK3+k3NWAJNZzxWcw4VD2n5xK8XKs1M
/894+4+xhhPZnoeAygmBq/zSW9B+Do1X/fAXbJSdzsWq0eiSCHL8WtsEVkpw
wBF/EpkqkQgQsN6UwOwyeOqYoh1lum+9feCPvVTtfkL+eOP6wVS1zBKc3E72
0X0hoZiZn7hXro0RwCR6rDnoiWYEtvhfuNjX9DlykwWjsC8ov3jXvf9JXGXF
NJwz422wbl3VeSbsvqS4shsBDHvCyBfi6EA6nwwTMEmUJ6jM1kXQRLE/RwXd
2/0VvLWtq5VA0QtgURovAMo0FimsVIjgc32u8Re7f/QahMqKuDz//NpO50tj
qrlqjEftLjjAudHJ1myfxPXg9cus6va2bVxisA0AefaaC4b78btC69chc4fC
IBF1DKwcoDMyVGnnpg66rCev4QAOprkViuNzBAitKKs1zA6lG3xzH3ytjy0v
0puxVk97E3jjOQNst0AJZ4ydR0hK2p7gISRM4oXnm0LvDG0A05wStQ8G+aDh
lRNC65Ci8iDzk6zqtEW2nRz1ZdJC0q4ky7jUVJ8HTmfU6Eyqn6y6gtnbVeaf
jGl8JL8bNKNxAXGRQFL0b5DD/mUhQWjh0LYvT0cSpRQT0bod0HjVF+YV7sRv
nont3IPkG6lfNOVKhUbpjiSXKNYd4O1Th8fSmMq7nrvqdl6zcytiAbxcymZt
DK0LvXY8extuzT2RSYq+FAHNuaONBlCuC851u4Tjq2WK/nHOirEAgqB+bFo0
YMONWy/hc5F3C/U5k8RUqJgUNTMkNScAvbCgCPsgSJna4KuYXLZEZYiiHEH+
jeaIzxZSyZHDKVx0IfoTPicNu5GfuWlAAjfgU0fvjqf+dP2hkk8Chm9DM9zE
E2jknheib2LJkHHXTo/HNZHOGKmdDhUB2TRPjhCYWh9jy1fivFHiCyeb1fHl
X0wB8yYyAqcbSYdfC2ckHez8b2iMg50mqy/t1iALYDfUskLZd9u0HOhQmMoi
oMqhzx4zSYjDJOXofi28t3tjEDFS/lv+j6ZWiy5/lcFU2XSbXREo7cLk75RF
0yf2TJXHv7jbeX5zN8XwTOUiERWthCSUMX+9mpg2/BZVPp8r+LoImdDmeAPd
qSXVuMQ1na3VNHKr83MY8wFPxfTNIqcXQiRNPLWwWXLnvyCNERD5Uttpgn/v
2G//OkYY1LxzRNNqoJzj4bsiYHdofEpOtY70zQor4DsJUo1SnldXmL58T/Gb
VHM9q++nLs30cXicYo7wdTLkclf+paWnjE2rB39gk9aU/FNJ3Xxsc6iVOKM4
UawBcumYh5dWBpz5ZBcFLpkDEckveTMv2MLbLsu8p1xrDre6omRZ8Q8dIn5x
F+jKnA2OZbXmVAmNn/CY3ddbEi08EkpgJW1CIbxcX+9q/VmVLDHYQSYLLe1N
f6R7kvVXwRN8MHN5EGtLNGBro5GadL+oW3cSbfzJbtgBKBZlnH1tBvyY7Aaz
YxHk15LYBiRqSHrL79dlq31uezKhK4h7TSs3ecCFqMzGj8oBpBfVvzJFep4U
aH2jIOL2QvlnsvdxzcG4Re57ljI7RNqFCZZVBWmYwTpnlhkT6skzF/lZP6OU
kPWtWpmgO0aUTlnIX62Dg3S14e5JqoGdWEQMHMV5nX5My22i0YMdlDZjGexh
jDalnlME1oLq8T7bA44KAewvtiSP+wAdiWcvsy9IeDO4UH8oE5uzk2qnsNeS
4kHTUbjwqVNkWU7sMkp2hV2fV+zxU1cqQnID8e00T8tT9kcSWvwb1Cd9a0t7
y9agdofZmsgn+ulaUtyGxFMXtawUUmQPCMRE3bdZPjJtawKwgbRnnh6TlYzi
uZZHpeK/enoNr4+ARGUL7XCgp+d4nyLGP4+TlXKGmBfbDwdL3jl6H2niMX1G
cCi474LvQQYHxVPd7KncVrxqONzgkVbHE1AQE6Ks4KCWKUQf5MrhYB3rqMYq
I5PW6DArsCi5tewHqtIN3qWIyFDdyPB9cDK1DVBpq1PrkUxffQtNROfJB5QB
V/W0jpsqle8W3P8abgEsAjClVArEmSbtYEWErX+Th/gwVeBaOO2791kiCIbU
4ZkV0RgW+///zZ7hsHAdMscNoCk8FtcIPPGD6nz6mnqRgXtY+lbuhCAnAhnH
SBmd9zY1dQqiUC+f7B+wkK4agChS7AKRZep35yByif8j/2+2UWzFod2rU+oZ
eiOZmiEKyk+YrRjN1VksHbJ8bwpbQNYkXxx4QHMrLq7mbGmGoMu0PFQGCJaT
K1yp279cJ8Gr0mcMFd7QbjSUQ3B1nItoG8dUEMjZBcOgMA7cm8SWV8R2KEBS
dGTABfqBgawMerkJRDwkaBGqQhsudF6dvxGAzPEzkZYrwNA2jXPx/mI64QH1
z2++Fs5LdxkR30U4+KtE/1LBEK2Hky4Y9V7YVsdJIau1U8SxYglOjMM+sSsu
Jrb0EOgxwbzpvHaGe4Vu2foxIZF7Ag1ydYOriFZphnZCZ9v0i6R6jWWYeUYs
l+dVybxkmX7R7BtDYSxxv3Cisx05q8ewFdq8yEP6AQ/uSmVl8YmocMuo8hxK
X+rq5QyILbHVzgh0ccbXGA8TSE17a2Id4GCmTFlKSBk1q1wCjENuul6WnFs6
TnKES1VWyXRiMwf9MqT6/T6rjH2s1Wm9vW9ZWLzxkZfY4bnN5mxHxFc38L5T
LF3f6cnEIJyNjc/JPHXAg2SgarLAEEVshG9Bej1c/7FNck1afgkkxN7Hh1YC
e68d2UScve5eXfTnckW+FZfhnqarT2/41hw0YfxsCR0CWzTny4alKMS/Fh52
q4y6hYd5Pb6ySOyJFiwOqLkIroJxdeu+chpoCrJTrKHmJ6ZWeEj0MJLeobKF
KywPORceMfL08hL4vb9NBS8bVOc7duGR3kMY34g4Uv75GN7egLdtFRNcpEMI
B1ycxf5K6dmgnp94W8x0acjWrIkuk5H9LUJZgx/hVWujwHQJcMz6ECSUMAaM
xzBYigWT7NWTb3FRP0CSPGNWEwdxSK631Odk3/iIuqaB+hJKERCgxgMKNgJq
a6gL7Ar+7tw9SIDkyYZNgHSArEUSQGjEwqriOKTHgADqPOUAAHD9uNBsxxtv
uekKcn657xgGQB1cOJ5jrXhri9sxCwb6Vhbnlj5PMJX5QCHlqO86fjod95mv
0xvLCNiauwx8CMZVY9ZM7eV7v4idWSdg5GmoL8jrvcCmAeDQYJbQB1I6bWrI
Cbc9ZAkVZgwlRJxuGtf9QXKEFnZOYHNgWEddNaRGlD4qvChvjJlHEIKHY/81
F1kc1aJFWabC2EeStX1/3QZsv4b6qFrCyfd08gxO+QV8ApGALYtPxZOGpfCC
RUOXBTcWu84qz25Iru//X1N31Kvo7PTGr0x4DdqQhksXA4M1btjN1p9ahyJe
002IH4KLFTri7TZGr5ZOsPk6iJYgK28FEB7lZeaQhXoitxHPb/yS9nOlHeX1
t+3VsJ8S4xYZlp+TWgpG/moLNN4Q7ahgdtYkB6/TxzTzlGRXOkLCCIuhIstL
DG6lTSXFwTIQLNMeC51FJ8636VaUH6zZGslooZ7To6IFkDnXmnt00bVOGThY
SQ3VqbKaKZt/uxU0IDFrFOz0SVJFEv7O9CCdsBb33f+VtIWtLrXtW7XXr3A7
UxPJb9Bb5W0aRbdFRxidUuPor5B1hWEAW02ZeaxOQVSs5vWKcETBLGdcPhCK
mVIUQfKOFlHHczgQp/Ge+oHBNGd7lM0CE2QFdGO4oeRRZdJMvk8GOHhqXkKC
S4kCg+hYDUqBu+D8cEI8OLR7jnlo4if1Dqsd5AWfsgLgZnB9797hI2tjqEj5
NO8TL43pgT8UQe5kUJQ1N5ezf5O+waILCe4urGviY6t6IpVGL+woQ140LULL
d3Qusze+YUriXVDoM9ttFDmUfse4d3Sbm4Yt//+FhGat7vrAMpaMFNtFDSrK
n41kfTBa5xcLhJTst360V3YRJF+ldOgTHI2RJmp/TgznfjOaLcI2IW1G4Dj5
UrlQAhWYOJd4ZhkedzsIwKlVt9r05pKf8voPRNveRCGlcJGEtdfr+74IgrBO
rFUWZhBchXXjTYBok493V9Y6CCjiRwYORJr4piyk1+J6vQbwgqTf+VrNXfBM
TgSDRmCd0y1+8V9SFFhjaUyvRkgUIWrhfi0Me2msMGKzcjFDGwRoJBMb82H0
rwoRkZggUqRKpvZlyTh9rEVSUzjj5LrzBltM3BJj2K5B91oupAXVY5s3Dc2m
zk++TsaCV0iEXg1xyMm+G8wPgHZrsS4p9hz4ZpGK3Prk9mq9osaZjaOAm4YJ
FaQJcMIWqmGwyzVTcyZ0vvgSAm2s37oRwdPF8QqhmL9cVGbeNz9Cj6f9bbDp
1tw3VYeUlvNs/QFWnPQ2RowXy2fYslanrzBDykqIyqcaJp7PWT6MIxCM6ZwY
nJ0LNSu9ZqawlvPNux3rb+KrwcTgjFzpe30+xcGCfy22WVQpXn3b/0S7FZEq
LJ7kq4chk1ZZjPteGlDhkSHurxbxPRxTX9kARjJ4DREIqBzqyfR9GBOyR5YB
GvW+5X7oDaozzP1E0XjEApBt8LM9QWxmySMcPrPo2Vi2fxy6tB2xwd7eAEVd
Hya3IPrSxuXHGAVtGkIn9XsTZ32PBJ8mNFsJDk4r+YIXJMnaDyaOjXBCXqvc
ZUNQV8XS6VFS9hwRHL9ZkeoVMAJwN13Zgy3CZsky218ydPp3N8uDvNECc4hE
KtaQvS0n12nYQOjfATWwh4dXQX7QZjaYegQ9kzmHqjlFcY+uujxb0JhpNeG5
4uY+ZwkBTN1YhgqxzPDhuJos9sFGZBpiqZoSceR6dSbhbehNIlX1LQU843w1
U/z/p7FPMuSv/Fr/B9/dyta9yd2DG+97aeprD+8KXyyxPvYLn9SSlGBImS4B
A6PRnlNtu6XtVcifkz87i0oFkan/N71hrDKmozIV0cvRRF+qT6rqXFFehGgz
PDqNGsaG+sohJGNbeKPRMoOq7LyE9f8/czYIUTwDEjwyoQRwU+arbtDs3HSz
o1YumOV4P/3OQcHAykc2TOfdvNjcuYW4A4kmhlaljvwsU2CBYtqWrDNv3D9t
gibdYP9qvb7CB3CpUx72E0fmZqixqzW3mGWKOm7BWizx6nFh3XfXdR2Y53HL
A7/vw1JdFZFzNdppHCM1ThNgl5RSuPoSYClNj5FsjdRHJ374SxWfdLzPj1tz
95uM6yVcU/WjIoBK3lW01nNgSeJsZVYvMBafCQOMF2RHjaespPKZn+CYOEt3
t5KoUTEYRbM1APoM5sR6TRwOseCaEeSoJZqvozndn+4ZkSEVwn3hDWFMCrGq
zxNm5bWsnlfNea3gELvoKDlsquit1VGaDWB8vBZwHkfULs3qn9zxXUhVUQB+
5drs3xTjEUHa1jmXsuMSnFNgCU1gVtjk/0upIy1LqyLeyqgMGCJRFAaQJBKV
C6WkSoc2+/WpLisYcy6pg4WbNrNuVz3610WgFHD2paFG9gjqJ0umUjgGyv7o
k5vt3V098/qhnH4i3s5ABkSouLf4ZKmyD9HPu6xqd9fcpUP2Yb2NTO78shnt
KkXa6Ur3Bfhfet/zHSHMcn83XZiXXLST9PIYyc01G3lj1qPr0AH67CeCjS3r
c2eE5quN5VEvSMg6ceAMw/SDf7QpJm2dC3n74TuDz51lOfiAAn/7OoyhgKSN
abaOcE4U+NTI/j67DdfOmjEmUS5HR2B1RXteldFHBbsygAsTruSOp0PuIJ+c
vqpi6mChd27Xa4c/1+ego7CfFvsZ/eaIkoXCFvCRiKJyadvlYPRHh0rv4hZX
jB8Iukj3aCC644P759b0p6f57Hwsrb3zj2mX2Dp2yBUb59lctH2VLMVqN9Fx
YD5olbRcnA0kR/oo1bSCfcp50Asoo3NABuPuzNIB3S0uaSRR21JXCZjlBS22
c7Ia/mpImMRUHUiYuIxfViI5bco+VLfmq/Arnmwl610A2FtyPATKmc7i8bt8
oLjAeHXLP/kVQPcQXRL63tOMKhwc3n+0TREmTi6vAJa8UpysHQuR8x+yMixz
Mc0z/TKtEQ6w3RWUInzuL3dLsGL0xNEtDV3UI6sW71gs5j6hIjkCYvzELeYy
DzJwtGxsj/LqrSVqxf6QfpcComuFeZCKWEOUP1a3XWn5B4z6Ozj/s/qIWjGe
EIJJ3Yngr2VpvuiWeQJe1617A1Uf4go8E1lHspSTvSSA5B0XJ56lW84KcaRY
psFwdNQE//Pdc2Ggc/JYmO5Z61sNpcn755reW/c5tSK2Cf/mAZs96xTcSpFA
eLyM+qes0A2vclHBiXqd6rxEe5kBVbzFZr3Eau8kLNJinUH+Uoh42GgTrrba
hqmp6mmJ4oB6RustNVOTjosWYOMFwJVeHdlfz3zXKKlnDDU6KvkI4XdFZlvJ
Gq4Q0GBn7LICb+1OYAkfHJSVcjZ6ITSSIQMUyUYE3YeESldUK3/fXaFLXeNP
NVGnM8DxCt8NutBBMRdNX8xuOnidSeXdRoBoJ5VdJtQ8QDuy7zqW0X/SGnia
z5x8rzxNd8IGK7vkg//7ly+3XXPYsmNI6gssRhvO/5/b8kNMLaivTenZRf0e
qVLOnCxdhOuc5ad7pxuQgelw+bFeZnyVUNh+LZsqplL1rTAR4AQCpttksFvi
HO9L7d5XPZmiLyip16MYsCW4Cf9d6t8Y087N2Jzacg22PVq2NM1+ZjMOx3I3
dXiICsx9iFow7wfjarkXX/GZ+d7s6F99FMHn9S82zNn0O7XNYP63L1/ORBR9
iU5XW/OligAXtPmyoJ6u0K4FV1vnb1+J/2iWI5Hg0zdcxkKzSW0s4R8i9aUQ
G8nybtoNe9GRyGyjtCTlEgHkS82BX5UVQaNPE9zqNCvXXKQ2Zi68HKQO46RZ
MJplepEb/tHroTjQyqVUq/pQVI2ILJ1RgnOZ8TDcLB8KYLnDF2B8UUjgX+22
13rn8CG6rA0pXcHC+ox6uQTP1hZai2eivt9qEZITP+w09WXeT4yesgzrCizy
v+Ib+4KFWV8DrXFYqqE6/XW50m4cdt3CLzD5hRd04aos2NZM7xGX7/uOxTxO
9oqrhJNYjDFdTnGUZ8RlqQ1kvT+EwS0iIuFdIgziYl63SDuGLzYD9gEQFAoD
ZAQp4nrE5XREEXmRQ4wRvwhnQKbSvoMIKEJjfb0I8oSNwhcr5Emmky6ZfjU6
tDL9lk3SnAPjVf9XPCDwKgqEzNmlpSf/uSNKULI+Phg6UzchqyEBjlXonVgm
efin204xjRgygWw0trHBX9kMs6CYREMmNZTi8ZqytuJ5f0943vfZqpxt+Wmq
7kYrSF7MxrftjGMim8D8+sfVWu7SWNeJ0Eqz9hU6K1HX70axn++KKhRcKGEf
hYiQU+VZT9r+uk97XCwDwtvMWmQwQl+D5hhRU4q0NPsTOHTOWhj6/ROHkCWV
s2sXoDsTWHijX15MNcLPsPeq6uJX1h3CmdWkh3SvKFIhCnHrlR7E6Gu9nTWj
Eu2Gh/7dlMBN7akcdtH3JlqikyA95CqBbvECRbi8epuTAtJYdfLsW1iwB6Ty
Pm1glorRUOt45tnLtsoJFFtNKcNNsgtNSBByYkXj+1KP7tp4u2AV7qrkAZWp
XYMLMuy421TskS6spjqamG8Xqoc3/XJcGwghehMoZlb+oC2RIP5wTupNC77K
5krpv/BEn9/Fh/BFeqdecMYwd3qWR2+UjNcOj/pPdM/R5iTWuSv02PwFpyao
g8YvGhIRUjkfPWcsa0WQoUdCj1PHX5+RZwlGUiXVB7r3Kiyi229mdXSW7xPf
oKmLhL0S17ZgKcJnc47ZEEaliWPjyKsdFp03aNOsA7FfiwkuMiqHAsrX9NIY
5PKCXK3bfYqPxpMxGcBEl3n9xgPcmaYDNMBcG5HWvRXiIc1pGRkPCPRmS7yR
EVWIH9gUfahshpZoIpRxlQWEKOxm4Oh0cPKTBNpIpFAmVlcRqRcb/FS/OI1m
SRuk1ikW8cQqgSUgiWjpTmLqHf8VGjZuVEqftVhUs/hJbPph6rSZpE/I7zwW
9BJS9A1rdiE6zuD6rOtXiz+iv/S6eZj1hrByc/087fKkAGAc+7xw6WmBC8xt
nHvqFXRaNA3FcnTpjw44a13FMbMBx/tTmJjPeXUCbD4j1j3aTwPeSgnmxTtg
sW5uamRVz3dx+MHNxecFHYlITWaJPkrornSl2eOk2xbdu2bKtgGxm9F0o2aE
ljzhkgjUvAXfSlFGwgCtGRP8MjxSw+oRW1oQU4JVVbAPoIjcyHfU3k93KtOe
bUceq3L+/FgUxiGYeLEg87Pi3T4bq1xqiO5XmiHs74t4OoLqaQ1rX/VGHz+u
lDL21rqZBXywxcbYt817e/lhPMcS+gMDMsov9f9mlwGV1gINw43YFwvGxqfr
HQz5cKzSUJz+0xzA7uLTcKc9s4njIf8QtRxfWPRu4psuzUmfcFM0CvFx6bgS
DVXWcNM1WBDGSOJA++MxiF1lUPt9RLG+aiWgLBN3mFlklV2r6cgMzUZKUD9D
QOhJmZXT9g0g2lD7/l71uKgdjgq7FehN9rMTiJMCXk2xnTJJ/0n5waG5TcSx
Jw7YmLnL+WztuhlgqnIrK6KtdMiveYQUxf1LM5Hid7LE4e8+Q0e7FjMeGgwi
wVqbWmBZiprdpP8QnozaAoIx/6vWjNuHfJ27WQM1jrPmeLPtxc6G6STiunNl
F1wgfH7qItQkuJZ5rXEE7q1r2fl07ZWVvhKCH3sqMKdHmjassJ8E9yjLi0/8
O1Ku52Co3DwX5kvxCS2tTwRh1zQkujWFs/z8e5xXdQp0AuEcfdjlBIeDKwGm
ttEsZLan+Vmxp0JIBSsakMSfval4oFyuNRuf4c1y6/1slyv3E3JuhlrywlBd
10Fc995BctX+pbuVym4MVljgOBc1awDAGLPALu7PwB4b/hG4Bxrj0PRkWPh2
kTs9tRhbz5nB4IdJpDtZ0WoOKm/0WVlM3Tob4vBAsaYImCdxb43HMkHhfthN
IzU+NJreDF9zzOyUQEjSovbxhX7f3pgW9zgf/+1QNUxQ7dy+N0lPClz86x4b
BykgzclDjjFvxckx0JITppIWkI7AI+hNcyZE5aoF8S3nVewqiGf/1Zbrieuc
tog1nmYc3yzzeHBcn2cnhJ1+xLEfXJGMqFf4XWEFfTEkNYFV4LQB1f7i6w2b
F69vd1O2IljqedjKi/10Dv+9fEbztFBJ6Y8o5P6YFZygapkOU88zczRG87jl
o1MHrG9CGVWKxmUsN+/UbuIPxXS4v0hZFOQ3O3GGsJtdtjGZDARb8XBLUqU3
AdfRvPsStWarTXnRYwCPSvt/INdQpvkWBQmwxaveEyUfne/TIdTOhJihniuj
ao3dkJa07dlwo21IgCRNHi6XgJh+vLy0YzKeb5psDSMib+T3eZeZ3MXlFkPW
n08Bmzbx/nG78YqyUih2PqJWdA9Nlx6NDm89blJFpdhBj9fWIYBZ204G9y2S
/xzK0UGlWE0z3VpaBAvMIeXxkN+WuNTT359wsP/OOlTrHWaFTDywMAulpTPK
vxfIdtrVOtv0XYefBEuPoIE17DrUXvfFDiyXojs+kv0H/5t9mfrVgzo9Xof1
8twCTWix892W/3TWWK1DZm+XqF1PNBt2htQWme+/JMnAKte2aMPm3edAHTof
cE4O/BrwvcAXPf5pFEQ5GQPSMXumL7sS2uOUL1IFCLhsxTnSsrGK9OXz/BzV
MIJtpx+UqCdUsMH2qe7AyGLgTRXpExexH20cZNJ88oxbZqffp3Yhuk9MZYLA
xaDwCLcG1ebx70lymRQMoegJC/5Qqc8tSxNLWXj2YHON7vSbC4afJygIIc7O
17oy6jZqp/PWGEZADSCUI0J6CrWszQsA9RoB9ZFGIcDTqk6M/0u9mkyA9Bdu
R5m307J9K7B4me0dhH/MONiOGBf5rLRmrsGN8K4hM07lH4nJsL5uhQnZo4Tw
Omj4YhGrIYhebHh1Expc+yZvO6s1Q3vpTjuFoj154RUzcUrcZD9VbTeTX4k4
TZOgySe1nFniewbOTpTGZL2CyWGcIExmpTmN82SJBCGqBm2HgklqPwSBp5sF
FwR7TqTu+4MNHQWoj6++0PYgrZN1Aqs1K03Dl3ikOlMRhXn6D5+J9LKCKuYX
rBRGrp0B6V5BHFBHN90GStFu80s69pywLWHKJ6OFEyzVs0sdyqcbgz4H7IX0
COZC/tQfVCINjAEc9dOc35Y9q+GyWyFU7uHrZUzdJZ9TSe30FuPGwIfGQ6zm
SnBy/ZpJQ3iS0JVvgBw80TToIEr26ADTtkg9G4h+Y+c8FKr9Gb9aTu/ulpqm
F4cbodL/Mt3yjxe0Lu/pXPYDiib6bO240pvxIaZRdK+V83faJWMKTIfMkdBz
nqz7drK8w8Lr1gKocTYuhxToDzHmW2rrbP9E3YaPwlpEEZMcnSAscVNcGd3B
EL2s4s+NNe10GX0njNuhthrOdDFqDP0OwjlHSzFP6yyjSYwEBQIpcsAd1OLh
lTBTcWm0ddOFBPXXG7oz8IwjOnHJ2qWpLy80AmLm0+R6Sz/55dXSCW0l47Y+
KooTNoJip9Me/+srKubUT73wT1PaGUvEo4+oWj3x+yWtHlF42YWXrk906gYF
DRvk0SjMkpdGp9qhgDCWIRLfs+yBFkgNQhmO4ZHIGeF0K69U2E88yNBhLSez
D5HaYBrYvMi56Klc/r1y5Uaavanai0l0ChcY3DlCDe/5xJ9NdHKk3yp6yf0i
u0ibtJ+9Glk+h53n9P4pQ6oc5TY9PH31SNccwTiEoRFK63HQc7biaGTCkuI6
a87/IE+8h/KtybCei2HoJhU9mK7UwJBUUhxSAxDbkI8otqifrstdWpUbOQ52
p7ftSkfSFf9RESAd36i5/8KpihD9xarQUOomhvDEygml3A7nMS1E1lZSh4SB
iC3JrUKcnT6QNZaNJQUU/H8kVkPbgyNoUK2AKN6tZlHU1VD1N48BhgIPQfO8
NZDkxuwPwqXlIrrby34aEglNGBfRc3bM0sJL2pmHhN97to5G2M4/C9GDioDp
k6Kgf/ZfxwxvGoUom5qyulh2zfnbH5dtcYBrPN0V2L+phZTp801oIYMxxmBh
wYlWMsqfSvUD5nrMOMQgowOYukaVTOx+kRRs1/pgLsHT/SDa56l7TQLLXyVt
5rYxlnrRSDYtOf+RCREq+sh5xUOb3YuB82b0Z9XHR+eIyupCHKiW2UHxSiql
YseZUxNZCUX53hVfVIiucWrgcPovpBlFVeDCUpanMdgKuu73g6hWEEMoZPLm
Or+jun9SS5CrkndqZekvMqMe1/mXiGfIS3gMgfOwg8oHO5mO+Ys6FdlKpdsF
CAl8Y8+vY1cz3rF7CoHpuLMe5uCdbhB5p4FuKQZr2cZW5aBnCQ+fnPJZ3m0R
xGX6JoBK0ZWkObRXrR7nxyBe8wn6TWZeKnS3QHmwY/xfxUrrM/kek4AemLp3
6Ud5s+GNOIyWE0jjYqIryJttgRrUBfWN+6x5vyjLVnPSWO5ykzuTVHB/Lkr7
3Vx40O2B/f0aHvY/m6DdVZ5o/eCv2AldvSCwt7l2iK4OSiMTZaJIvOtEI4pX
s24YlwQiZalLA7geOxpQOT4ZVxSPXMTOy/XNHXJ9Hk2fZgLwTIjPTsCVHgmI
2jKm7ep/1mrSAdUS2HdV3BZ/U16JWWJI54Xbg+GWQQbRbrp422B6IP5m4G9g
RkJ5gFt2nPUGtSpPd6TRzSDtq3czuy9MEDeOsa1Kq3RWiLgiS+dgEYnZQ1HK
9bc3apaxQt8TtUuoYl3vF4JVMjp4DNn3H98QWiiZQ/d4knddxEzWgKPcTRPX
H4ZwKt/xOEjrQCYEFemQX4uDhg0x8JsKUEzE+opQSsPOiGOi7ASgCcO37DHa
59UAM95B/SlIn7IoFCcbfUl3EV6oIKWDNerE2/rJrApVThL04Q+3yxcPJJo7
eTQZn+qrDDi1yWomNe6fPiG2DW0780VTZreuzInk9LdO1s1FX2KA2c2Pf4tz
vX/Gop4U8hzi4yKDwWF+MQYo4/DKF/t1Cz5pS0sRgLBNFv0=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "OJXsOzX3SCOyhcBXS9yryN9cWQxQkhDHUr4mzQikLKNKnB6JkSYY9xNnmYkvVOJ5f3SnsxLM71tWjwpqmyTCVkTt4jikDmXDCnl6lQn2TVy78ivgbebFE/F7GUr3Z8AASPmtz4v12cD/Cz7nTJMTG81IGzEoV1S4KsV3MBcbB+1TqTshtjzQ4oMMPpNw9ltjOjjqx8CktvtqLiQWjnKfQh8i3R/5yQlzObBDq+VCqAPsTnYdflrq4Ab4rxhnHhTDx1MBCTvCpkDVWd7rNwq7cljRgMrF9H4gnHVaV6EdSViy2cmnFEUDMtY27uzFc2okvb3RRMH8QjnW0vKMbPSZwKmVRxjbHO8AOrFGcKxKaK4iGGoE7rzhKjDloW6TbdtGA4D+Q2e0yG4OelzERF/Kwkce1Ctu16NiB8gUhf/mjyO9IShvvSLzsQ7yuUhdxCA2mXYPrnyRIajzyVXywrPAfrUFB0C63iMkW99OurQo7/NXUOLC+pC2j2CFWrU+xp/AqkHpPa6wox6idOtjbSHDb7ljFFQ2CJaQk4T7pfVOeF02e8hScftK8gxD9SryRI+Hb5pckk/W/+zpdtzPbVJdB6wRk5UefATWJhqhDcqmIksdQRlnBsKdXX+dzNosqfHri5uNxUMMgpB1IEk88LkFVMw6ScnDDhwL98+pwgPTwiS6CfQmzevSDTJeqWKOTemG6NzKEEfMLyRp24SizkocXIp5BN1HuwmHz7ggFvPL+qjjBfy4iDnaxaH+QpHm7OEXvnSBxUGGD7pDTqBgAd3Lv88cBS0/ppzY4eH7SazFd2SpV4rZzCShgd/6ZT0NyQXq6wlIba677IEd+twTyM8t3FLpzoNKZdplBBZGsY8N6oClA8tmoZ1GqqJE7ENrD3TDgVGJAF14OT+8/+jZvSPjmYQyzPQHvwqyp+1WOh4xkGPDAhplAyjFJNQxgJ6Mj1BnfZMka6q1kTBg79RW8Kwuqpf1D9jPR3KTpQM6iFhbO6ltFmLRRR0xSHSh21uE9AW8"
`endif